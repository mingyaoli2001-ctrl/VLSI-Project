* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : MAC                                          *
* Netlisted  : Sat Dec 13 12:39:58 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765647593020                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765647593020 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765647593020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765647593021                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765647593021 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765647593021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765647593022                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765647593022 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765647593022

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765647593023                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765647593023 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765647593023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765647593024                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765647593024 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765647593024

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765647593025                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765647593025 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765647593025

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765647593026                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765647593026 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765647593026

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765647593027                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765647593027 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765647593027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765647593028                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765647593028 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765647593028

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765647593029                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765647593029 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765647593029

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930210                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930210 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930211                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930211 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930211

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930212                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930212 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930212

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656475930214                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656475930214 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656475930214

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656475930215                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656475930215 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656475930215

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930216                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930216 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930216

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765647593020                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765647593020 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765647593020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593021                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593021 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X0 4 M3_M2_CDNS_765647593026 $T=1850 2810 0 90 $X=1600 $Y=2590
X1 4 M4_M3_CDNS_765647593027 $T=1850 2810 0 90 $X=1600 $Y=2590
X2 4 M5_M4_CDNS_765647593028 $T=1850 2810 0 90 $X=1600 $Y=2590
X3 4 M6_M5_CDNS_765647593029 $T=1850 2810 0 90 $X=1600 $Y=2590
X4 4 M2_M1_CDNS_7656475930210 $T=1850 2810 0 90 $X=1600 $Y=2590
X5 6 M2_M1_CDNS_7656475930211 $T=690 3330 0 0 $X=610 $Y=3200
X6 1 M2_M1_CDNS_7656475930211 $T=1190 1490 0 0 $X=1110 $Y=1360
X7 1 M2_M1_CDNS_7656475930211 $T=2520 1490 0 0 $X=2440 $Y=1360
X8 6 M2_M1_CDNS_7656475930211 $T=2550 3330 0 0 $X=2470 $Y=3200
X9 1 M1_PO_CDNS_7656475930214 $T=320 1490 0 0 $X=220 $Y=1240
X10 5 M1_PO_CDNS_7656475930214 $T=1540 2050 0 0 $X=1440 $Y=1800
X11 5 M1_PO_CDNS_7656475930214 $T=3400 2050 0 0 $X=3300 $Y=1800
X12 7 M1_PO_CDNS_7656475930215 $T=2470 2570 0 0 $X=2370 $Y=2450
X13 1 M2_M1_CDNS_7656475930216 $T=320 1490 0 0 $X=240 $Y=1240
X14 5 M2_M1_CDNS_7656475930216 $T=1540 2050 0 0 $X=1460 $Y=1800
X15 5 M2_M1_CDNS_7656475930216 $T=3400 2050 0 0 $X=3320 $Y=1800
X16 2 2 1 6 3 pmos1v_CDNS_765647593020 $T=420 3660 0 0 $X=0 $Y=3460
X17 1 2 5 4 3 pmos1v_CDNS_765647593020 $T=1350 3660 0 0 $X=930 $Y=3460
X18 6 2 7 4 3 pmos1v_CDNS_765647593020 $T=2370 3660 1 180 $X=1860 $Y=3460
X19 2 2 5 7 3 pmos1v_CDNS_765647593020 $T=3300 3660 1 180 $X=2790 $Y=3460
X20 3 3 1 6 nmos1v_CDNS_765647593021 $T=420 800 0 0 $X=0 $Y=240
X21 4 3 5 6 nmos1v_CDNS_765647593021 $T=1440 800 1 180 $X=930 $Y=240
X22 4 3 7 1 nmos1v_CDNS_765647593021 $T=2280 800 0 0 $X=1860 $Y=240
X23 3 3 5 7 nmos1v_CDNS_765647593021 $T=3300 800 1 180 $X=2790 $Y=240
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656475930217                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656475930217 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656475930217

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930218                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930218 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930218

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593022                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593022 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593022

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765647593023                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765647593023 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765647593023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593024                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593024 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593024

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765647593025                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765647593025 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765647593025

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765647593026                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765647593026 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765647593026

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593027                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593027 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=3
X0 1 M2_M1_CDNS_7656475930211 $T=1510 -2070 0 0 $X=1430 $Y=-2200
X1 1 M2_M1_CDNS_7656475930211 $T=3010 -2070 0 0 $X=2930 $Y=-2200
X2 2 M1_PO_CDNS_7656475930215 $T=1870 -1670 0 0 $X=1770 $Y=-1790
X3 1 M1_PO_CDNS_7656475930215 $T=2510 -2070 0 0 $X=2410 $Y=-2190
X4 6 M1_PO_CDNS_7656475930215 $T=4500 -2020 0 0 $X=4400 $Y=-2140
X5 5 M3_M2_CDNS_7656475930217 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X6 5 M2_M1_CDNS_7656475930218 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X7 4 5 6 nmos1v_CDNS_765647593022 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X8 3 5 6 4 pmos1v_CDNS_765647593023 $T=4560 -1510 0 0 $X=3880 $Y=-1710
X9 4 1 7 nmos1v_CDNS_765647593024 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X10 3 2 6 4 pmos1v_CDNS_765647593025 $T=1930 -1320 0 0 $X=1250 $Y=-1520
X11 3 6 1 4 pmos1v_CDNS_765647593026 $T=2430 -1320 1 180 $X=1980 $Y=-1520
X12 6 2 7 4 nmos1v_CDNS_765647593027 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656475930219                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656475930219 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656475930219

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656475930220                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656475930220 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656475930220

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656475930221                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656475930221 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656475930221

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656475930222                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656475930222 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656475930222

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656475930223                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656475930223 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656475930223

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656475930224                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656475930224 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656475930224

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930226                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930226 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930226

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656475930227                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656475930227 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656475930227

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656475930228                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656475930228 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656475930228

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656475930229                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656475930229 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656475930229

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656475930230                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656475930230 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656475930230

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656475930231                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656475930231 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656475930231

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765647593028                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765647593028 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 4 3 1 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765647593028

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593029                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593029 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593029

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39
*.DEVICECLIMB
** N=39 EP=39 FDC=54
X0 2 M3_M2_CDNS_765647593020 $T=610 4030 0 0 $X=530 $Y=3780
X1 1 M3_M2_CDNS_765647593020 $T=930 5440 0 0 $X=850 $Y=5190
X2 2 M3_M2_CDNS_765647593020 $T=2790 4030 0 0 $X=2710 $Y=3780
X3 7 M3_M2_CDNS_765647593020 $T=3110 3560 0 0 $X=3030 $Y=3310
X4 8 M3_M2_CDNS_765647593020 $T=4110 1490 0 0 $X=4030 $Y=1240
X5 1 M3_M2_CDNS_765647593020 $T=5580 5440 0 0 $X=5500 $Y=5190
X6 2 M3_M2_CDNS_765647593020 $T=7440 4030 0 0 $X=7360 $Y=3780
X7 10 M3_M2_CDNS_765647593020 $T=8700 3090 0 0 $X=8620 $Y=2840
X8 11 M3_M2_CDNS_765647593020 $T=9690 1490 0 0 $X=9610 $Y=1240
X9 9 M3_M2_CDNS_765647593020 $T=10230 6380 0 0 $X=10150 $Y=6130
X10 1 M3_M2_CDNS_765647593020 $T=12090 5440 0 0 $X=12010 $Y=5190
X11 2 M3_M2_CDNS_765647593020 $T=13950 4030 0 0 $X=13870 $Y=3780
X12 10 M3_M2_CDNS_765647593020 $T=15810 3090 0 0 $X=15730 $Y=2840
X13 13 M3_M2_CDNS_765647593020 $T=17130 1490 0 0 $X=17050 $Y=1240
X14 14 M3_M2_CDNS_765647593020 $T=17490 2630 0 0 $X=17410 $Y=2380
X15 9 M3_M2_CDNS_765647593020 $T=18600 6380 0 0 $X=18520 $Y=6130
X16 1 M3_M2_CDNS_765647593020 $T=20460 5440 0 0 $X=20380 $Y=5190
X17 2 M3_M2_CDNS_765647593020 $T=22320 4030 0 0 $X=22240 $Y=3780
X18 10 M3_M2_CDNS_765647593020 $T=24180 3090 0 0 $X=24100 $Y=2840
X19 15 M3_M2_CDNS_765647593020 $T=26430 1490 0 0 $X=26350 $Y=1240
X20 2 M4_M3_CDNS_765647593021 $T=610 4030 0 0 $X=530 $Y=3780
X21 1 M4_M3_CDNS_765647593021 $T=930 5440 0 0 $X=850 $Y=5190
X22 2 M4_M3_CDNS_765647593021 $T=2790 4030 0 0 $X=2710 $Y=3780
X23 1 M4_M3_CDNS_765647593021 $T=5580 5440 0 0 $X=5500 $Y=5190
X24 2 M4_M3_CDNS_765647593021 $T=7440 4030 0 0 $X=7360 $Y=3780
X25 10 M4_M3_CDNS_765647593021 $T=8700 3090 0 0 $X=8620 $Y=2840
X26 9 M4_M3_CDNS_765647593021 $T=10230 6380 0 0 $X=10150 $Y=6130
X27 1 M4_M3_CDNS_765647593021 $T=12090 5440 0 0 $X=12010 $Y=5190
X28 2 M4_M3_CDNS_765647593021 $T=13950 4030 0 0 $X=13870 $Y=3780
X29 10 M4_M3_CDNS_765647593021 $T=15810 3090 0 0 $X=15730 $Y=2840
X30 9 M4_M3_CDNS_765647593021 $T=18600 6380 0 0 $X=18520 $Y=6130
X31 1 M4_M3_CDNS_765647593021 $T=20460 5440 0 0 $X=20380 $Y=5190
X32 2 M4_M3_CDNS_765647593021 $T=22320 4030 0 0 $X=22240 $Y=3780
X33 10 M4_M3_CDNS_765647593021 $T=24180 3090 0 0 $X=24100 $Y=2840
X34 7 M4_M3_CDNS_765647593025 $T=3110 3560 0 0 $X=3030 $Y=3310
X35 8 M4_M3_CDNS_765647593025 $T=4110 1490 0 0 $X=4030 $Y=1240
X36 11 M4_M3_CDNS_765647593025 $T=9690 1490 0 0 $X=9610 $Y=1240
X37 13 M4_M3_CDNS_765647593025 $T=17130 1490 0 0 $X=17050 $Y=1240
X38 14 M4_M3_CDNS_765647593025 $T=17490 2630 0 0 $X=17410 $Y=2380
X39 15 M4_M3_CDNS_765647593025 $T=26430 1490 0 0 $X=26350 $Y=1240
X40 16 M3_M2_CDNS_765647593026 $T=3580 4500 0 0 $X=3360 $Y=4250
X41 17 M3_M2_CDNS_765647593026 $T=9160 4500 0 0 $X=8940 $Y=4250
X42 18 M3_M2_CDNS_765647593026 $T=16600 4500 0 0 $X=16380 $Y=4250
X43 19 M3_M2_CDNS_765647593026 $T=25900 4500 0 0 $X=25680 $Y=4250
X44 16 M4_M3_CDNS_765647593027 $T=3580 4500 0 0 $X=3360 $Y=4250
X45 17 M4_M3_CDNS_765647593027 $T=9160 4500 0 0 $X=8940 $Y=4250
X46 18 M4_M3_CDNS_765647593027 $T=16600 4500 0 0 $X=16380 $Y=4250
X47 19 M4_M3_CDNS_765647593027 $T=25900 4500 0 0 $X=25680 $Y=4250
X48 16 M5_M4_CDNS_765647593028 $T=3580 4500 0 0 $X=3360 $Y=4250
X49 17 M5_M4_CDNS_765647593028 $T=9160 4500 0 0 $X=8940 $Y=4250
X50 18 M5_M4_CDNS_765647593028 $T=16600 4500 0 0 $X=16380 $Y=4250
X51 19 M5_M4_CDNS_765647593028 $T=25900 4500 0 0 $X=25680 $Y=4250
X52 16 M2_M1_CDNS_7656475930210 $T=3580 4500 0 0 $X=3360 $Y=4250
X53 17 M2_M1_CDNS_7656475930210 $T=9160 4500 0 0 $X=8940 $Y=4250
X54 18 M2_M1_CDNS_7656475930210 $T=16600 4500 0 0 $X=16380 $Y=4250
X55 19 M2_M1_CDNS_7656475930210 $T=25900 4500 0 0 $X=25680 $Y=4250
X56 2 M2_M1_CDNS_7656475930212 $T=610 4030 0 0 $X=530 $Y=3780
X57 1 M2_M1_CDNS_7656475930212 $T=930 5440 0 0 $X=850 $Y=5190
X58 3 M2_M1_CDNS_7656475930212 $T=1860 4970 0 0 $X=1780 $Y=4720
X59 2 M2_M1_CDNS_7656475930212 $T=2790 4030 0 0 $X=2710 $Y=3780
X60 7 M2_M1_CDNS_7656475930212 $T=3110 3560 0 0 $X=3030 $Y=3310
X61 8 M2_M1_CDNS_7656475930212 $T=4110 1490 0 0 $X=4030 $Y=1240
X62 6 M2_M1_CDNS_7656475930212 $T=4650 5910 0 0 $X=4570 $Y=5660
X63 1 M2_M1_CDNS_7656475930212 $T=5580 5440 0 0 $X=5500 $Y=5190
X64 3 M2_M1_CDNS_7656475930212 $T=6510 4970 0 0 $X=6430 $Y=4720
X65 2 M2_M1_CDNS_7656475930212 $T=7440 4030 0 0 $X=7360 $Y=3780
X66 7 M2_M1_CDNS_7656475930212 $T=8370 3560 0 0 $X=8290 $Y=3310
X67 10 M2_M1_CDNS_7656475930212 $T=8700 3090 0 0 $X=8620 $Y=2840
X68 11 M2_M1_CDNS_7656475930212 $T=9690 1490 0 0 $X=9610 $Y=1240
X69 9 M2_M1_CDNS_7656475930212 $T=10230 6380 0 0 $X=10150 $Y=6130
X70 6 M2_M1_CDNS_7656475930212 $T=11160 5910 0 0 $X=11080 $Y=5660
X71 1 M2_M1_CDNS_7656475930212 $T=12090 5440 0 0 $X=12010 $Y=5190
X72 3 M2_M1_CDNS_7656475930212 $T=13020 4970 0 0 $X=12940 $Y=4720
X73 2 M2_M1_CDNS_7656475930212 $T=13950 4030 0 0 $X=13870 $Y=3780
X74 7 M2_M1_CDNS_7656475930212 $T=14880 3560 0 0 $X=14800 $Y=3310
X75 10 M2_M1_CDNS_7656475930212 $T=15810 3090 0 0 $X=15730 $Y=2840
X76 13 M2_M1_CDNS_7656475930212 $T=17130 1490 0 0 $X=17050 $Y=1240
X77 14 M2_M1_CDNS_7656475930212 $T=17490 2630 0 0 $X=17410 $Y=2380
X78 12 M2_M1_CDNS_7656475930212 $T=17670 6850 0 0 $X=17590 $Y=6600
X79 9 M2_M1_CDNS_7656475930212 $T=18600 6380 0 0 $X=18520 $Y=6130
X80 6 M2_M1_CDNS_7656475930212 $T=19530 5910 0 0 $X=19450 $Y=5660
X81 1 M2_M1_CDNS_7656475930212 $T=20460 5440 0 0 $X=20380 $Y=5190
X82 3 M2_M1_CDNS_7656475930212 $T=21390 4970 0 0 $X=21310 $Y=4720
X83 2 M2_M1_CDNS_7656475930212 $T=22320 4030 0 0 $X=22240 $Y=3780
X84 7 M2_M1_CDNS_7656475930212 $T=23250 3560 0 0 $X=23170 $Y=3310
X85 10 M2_M1_CDNS_7656475930212 $T=24180 3090 0 0 $X=24100 $Y=2840
X86 14 M2_M1_CDNS_7656475930212 $T=25110 2620 0 0 $X=25030 $Y=2370
X87 15 M2_M1_CDNS_7656475930212 $T=26430 1490 0 0 $X=26350 $Y=1240
X88 4 4 2 20 5 pmos1v_CDNS_765647593020 $T=2980 8370 1 180 $X=2470 $Y=8170
X89 4 4 16 8 5 pmos1v_CDNS_765647593020 $T=3820 8370 0 0 $X=3400 $Y=8170
X90 4 4 6 17 5 pmos1v_CDNS_765647593020 $T=4750 8370 0 0 $X=4330 $Y=8170
X91 21 4 3 17 5 pmos1v_CDNS_765647593020 $T=6700 8370 1 180 $X=6190 $Y=8170
X92 22 4 2 21 5 pmos1v_CDNS_765647593020 $T=7630 8370 1 180 $X=7120 $Y=8170
X93 4 4 7 22 5 pmos1v_CDNS_765647593020 $T=8560 8370 1 180 $X=8050 $Y=8170
X94 4 4 17 11 5 pmos1v_CDNS_765647593020 $T=9400 8370 0 0 $X=8980 $Y=8170
X95 4 4 9 18 5 pmos1v_CDNS_765647593020 $T=10330 8370 0 0 $X=9910 $Y=8170
X96 23 4 6 18 5 pmos1v_CDNS_765647593020 $T=11350 8370 1 180 $X=10840 $Y=8170
X97 24 4 1 18 5 pmos1v_CDNS_765647593020 $T=12280 8370 1 180 $X=11770 $Y=8170
X98 25 4 3 18 5 pmos1v_CDNS_765647593020 $T=13210 8370 1 180 $X=12700 $Y=8170
X99 24 4 2 25 5 pmos1v_CDNS_765647593020 $T=14140 8370 1 180 $X=13630 $Y=8170
X100 23 4 7 24 5 pmos1v_CDNS_765647593020 $T=15070 8370 1 180 $X=14560 $Y=8170
X101 4 4 10 23 5 pmos1v_CDNS_765647593020 $T=16000 8370 1 180 $X=15490 $Y=8170
X102 4 4 12 19 5 pmos1v_CDNS_765647593020 $T=17770 8370 0 0 $X=17350 $Y=8170
X103 26 4 6 19 5 pmos1v_CDNS_765647593020 $T=19720 8370 1 180 $X=19210 $Y=8170
X104 27 4 1 19 5 pmos1v_CDNS_765647593020 $T=20650 8370 1 180 $X=20140 $Y=8170
X105 27 4 2 28 5 pmos1v_CDNS_765647593020 $T=22510 8370 1 180 $X=22000 $Y=8170
X106 26 4 7 27 5 pmos1v_CDNS_765647593020 $T=23440 8370 1 180 $X=22930 $Y=8170
X107 4 4 14 29 5 pmos1v_CDNS_765647593020 $T=25300 8370 1 180 $X=24790 $Y=8170
X108 4 4 19 15 5 pmos1v_CDNS_765647593020 $T=26140 8370 0 0 $X=25720 $Y=8170
X109 5 5 1 30 nmos1v_CDNS_765647593021 $T=1030 800 0 0 $X=610 $Y=240
X110 30 5 3 16 nmos1v_CDNS_765647593021 $T=1960 800 0 0 $X=1540 $Y=240
X111 5 5 6 31 nmos1v_CDNS_765647593021 $T=4750 800 0 0 $X=4330 $Y=240
X112 31 5 2 17 nmos1v_CDNS_765647593021 $T=7540 800 0 0 $X=7120 $Y=240
X113 5 5 7 17 nmos1v_CDNS_765647593021 $T=8560 800 1 180 $X=8050 $Y=240
X114 5 5 17 11 nmos1v_CDNS_765647593021 $T=9400 800 0 0 $X=8980 $Y=240
X115 32 5 1 33 nmos1v_CDNS_765647593021 $T=12190 800 0 0 $X=11770 $Y=240
X116 33 5 3 18 nmos1v_CDNS_765647593021 $T=13120 800 0 0 $X=12700 $Y=240
X117 34 5 7 18 nmos1v_CDNS_765647593021 $T=14980 800 0 0 $X=14560 $Y=240
X118 5 5 10 18 nmos1v_CDNS_765647593021 $T=16000 800 1 180 $X=15490 $Y=240
X119 5 5 18 13 nmos1v_CDNS_765647593021 $T=16840 800 0 0 $X=16420 $Y=240
X120 35 5 9 36 nmos1v_CDNS_765647593021 $T=18700 800 0 0 $X=18280 $Y=240
X121 36 5 7 19 nmos1v_CDNS_765647593021 $T=23350 800 0 0 $X=22930 $Y=240
X122 5 5 19 15 nmos1v_CDNS_765647593021 $T=26140 800 0 0 $X=25720 $Y=240
X123 3 M3_M2_CDNS_7656475930217 $T=250 4970 0 90 $X=0 $Y=4890
X124 3 M3_M2_CDNS_7656475930217 $T=1860 4970 0 0 $X=1780 $Y=4720
X125 6 M3_M2_CDNS_7656475930217 $T=4650 5910 0 0 $X=4570 $Y=5660
X126 3 M3_M2_CDNS_7656475930217 $T=6510 4970 0 0 $X=6430 $Y=4720
X127 7 M3_M2_CDNS_7656475930217 $T=8370 3560 0 0 $X=8290 $Y=3310
X128 6 M3_M2_CDNS_7656475930217 $T=11160 5910 0 0 $X=11080 $Y=5660
X129 3 M3_M2_CDNS_7656475930217 $T=13020 4970 0 0 $X=12940 $Y=4720
X130 7 M3_M2_CDNS_7656475930217 $T=14880 3560 0 0 $X=14800 $Y=3310
X131 12 M3_M2_CDNS_7656475930217 $T=17670 6850 0 0 $X=17590 $Y=6600
X132 6 M3_M2_CDNS_7656475930217 $T=19530 5910 0 0 $X=19450 $Y=5660
X133 3 M3_M2_CDNS_7656475930217 $T=21390 4970 0 0 $X=21310 $Y=4720
X134 7 M3_M2_CDNS_7656475930217 $T=23250 3560 0 0 $X=23170 $Y=3310
X135 14 M3_M2_CDNS_7656475930217 $T=25110 2620 0 0 $X=25030 $Y=2370
X136 3 M2_M1_CDNS_7656475930218 $T=250 4970 0 90 $X=0 $Y=4890
X137 1 M4_M3_CDNS_7656475930219 $T=80 5580 0 0 $X=0 $Y=5190
X138 16 M4_M3_CDNS_7656475930219 $T=1540 7840 0 0 $X=1460 $Y=7450
X139 6 M4_M3_CDNS_7656475930219 $T=2130 6050 0 0 $X=2050 $Y=5660
X140 16 M4_M3_CDNS_7656475930219 $T=2470 1570 0 0 $X=2390 $Y=1180
X141 17 M4_M3_CDNS_7656475930219 $T=5260 7840 0 0 $X=5180 $Y=7450
X142 17 M4_M3_CDNS_7656475930219 $T=6450 7840 0 0 $X=6370 $Y=7450
X143 17 M4_M3_CDNS_7656475930219 $T=6860 1570 0 0 $X=6780 $Y=1180
X144 9 M4_M3_CDNS_7656475930219 $T=7710 6520 0 0 $X=7630 $Y=6130
X145 17 M4_M3_CDNS_7656475930219 $T=8050 1570 0 0 $X=7970 $Y=1180
X146 18 M4_M3_CDNS_7656475930219 $T=10840 7840 0 0 $X=10760 $Y=7450
X147 18 M4_M3_CDNS_7656475930219 $T=12030 7840 0 0 $X=11950 $Y=7450
X148 18 M4_M3_CDNS_7656475930219 $T=12960 7840 0 0 $X=12880 $Y=7450
X149 18 M4_M3_CDNS_7656475930219 $T=13370 1570 0 0 $X=13290 $Y=1180
X150 18 M4_M3_CDNS_7656475930219 $T=14300 1570 0 0 $X=14220 $Y=1180
X151 18 M4_M3_CDNS_7656475930219 $T=15490 1570 0 0 $X=15410 $Y=1180
X152 12 M4_M3_CDNS_7656475930219 $T=16080 6990 0 0 $X=16000 $Y=6600
X153 19 M4_M3_CDNS_7656475930219 $T=18280 7840 0 0 $X=18200 $Y=7450
X154 19 M4_M3_CDNS_7656475930219 $T=19470 7840 0 0 $X=19390 $Y=7450
X155 19 M4_M3_CDNS_7656475930219 $T=20400 7840 0 0 $X=20320 $Y=7450
X156 19 M4_M3_CDNS_7656475930219 $T=21330 7840 0 0 $X=21250 $Y=7450
X157 19 M4_M3_CDNS_7656475930219 $T=21740 1570 0 0 $X=21660 $Y=1180
X158 19 M4_M3_CDNS_7656475930219 $T=22670 1570 0 0 $X=22590 $Y=1180
X159 19 M4_M3_CDNS_7656475930219 $T=23600 1570 0 0 $X=23520 $Y=1180
X160 19 M4_M3_CDNS_7656475930219 $T=24790 1570 0 0 $X=24710 $Y=1180
X161 16 M7_M6_CDNS_7656475930220 $T=1540 7840 0 0 $X=1460 $Y=7450
X162 16 M7_M6_CDNS_7656475930220 $T=2470 1570 0 0 $X=2390 $Y=1180
X163 17 M7_M6_CDNS_7656475930220 $T=5260 7840 0 0 $X=5180 $Y=7450
X164 17 M7_M6_CDNS_7656475930220 $T=6450 7840 0 0 $X=6370 $Y=7450
X165 17 M7_M6_CDNS_7656475930220 $T=6860 1570 0 0 $X=6780 $Y=1180
X166 17 M7_M6_CDNS_7656475930220 $T=8050 1570 0 0 $X=7970 $Y=1180
X167 18 M7_M6_CDNS_7656475930220 $T=10840 7840 0 0 $X=10760 $Y=7450
X168 18 M7_M6_CDNS_7656475930220 $T=12030 7840 0 0 $X=11950 $Y=7450
X169 18 M7_M6_CDNS_7656475930220 $T=12960 7840 0 0 $X=12880 $Y=7450
X170 18 M7_M6_CDNS_7656475930220 $T=13370 1570 0 0 $X=13290 $Y=1180
X171 18 M7_M6_CDNS_7656475930220 $T=14300 1570 0 0 $X=14220 $Y=1180
X172 18 M7_M6_CDNS_7656475930220 $T=15490 1570 0 0 $X=15410 $Y=1180
X173 19 M7_M6_CDNS_7656475930220 $T=18280 7840 0 0 $X=18200 $Y=7450
X174 19 M7_M6_CDNS_7656475930220 $T=19470 7840 0 0 $X=19390 $Y=7450
X175 19 M7_M6_CDNS_7656475930220 $T=20400 7840 0 0 $X=20320 $Y=7450
X176 19 M7_M6_CDNS_7656475930220 $T=21330 7840 0 0 $X=21250 $Y=7450
X177 19 M7_M6_CDNS_7656475930220 $T=21740 1570 0 0 $X=21660 $Y=1180
X178 19 M7_M6_CDNS_7656475930220 $T=22670 1570 0 0 $X=22590 $Y=1180
X179 19 M7_M6_CDNS_7656475930220 $T=23600 1570 0 0 $X=23520 $Y=1180
X180 19 M7_M6_CDNS_7656475930220 $T=24790 1570 0 0 $X=24710 $Y=1180
X181 16 M1_PO_CDNS_7656475930221 $T=3580 4500 0 0 $X=3340 $Y=4250
X182 17 M1_PO_CDNS_7656475930221 $T=9160 4500 0 0 $X=8920 $Y=4250
X183 18 M1_PO_CDNS_7656475930221 $T=16600 4500 0 0 $X=16360 $Y=4250
X184 16 M6_M5_CDNS_7656475930222 $T=3580 4500 0 0 $X=3360 $Y=4250
X185 17 M6_M5_CDNS_7656475930222 $T=9160 4500 0 0 $X=8940 $Y=4250
X186 18 M6_M5_CDNS_7656475930222 $T=16600 4500 0 0 $X=16380 $Y=4250
X187 19 M6_M5_CDNS_7656475930222 $T=25900 4500 0 0 $X=25680 $Y=4250
X188 2 M5_M4_CDNS_7656475930223 $T=610 4030 0 0 $X=530 $Y=3780
X189 1 M5_M4_CDNS_7656475930223 $T=930 5440 0 0 $X=850 $Y=5190
X190 2 M5_M4_CDNS_7656475930223 $T=2790 4030 0 0 $X=2710 $Y=3780
X191 1 M5_M4_CDNS_7656475930223 $T=5580 5440 0 0 $X=5500 $Y=5190
X192 2 M5_M4_CDNS_7656475930223 $T=7440 4030 0 0 $X=7360 $Y=3780
X193 10 M5_M4_CDNS_7656475930223 $T=8700 3090 0 0 $X=8620 $Y=2840
X194 9 M5_M4_CDNS_7656475930223 $T=10230 6380 0 0 $X=10150 $Y=6130
X195 1 M5_M4_CDNS_7656475930223 $T=12090 5440 0 0 $X=12010 $Y=5190
X196 2 M5_M4_CDNS_7656475930223 $T=13950 4030 0 0 $X=13870 $Y=3780
X197 10 M5_M4_CDNS_7656475930223 $T=15810 3090 0 0 $X=15730 $Y=2840
X198 9 M5_M4_CDNS_7656475930223 $T=18600 6380 0 0 $X=18520 $Y=6130
X199 1 M5_M4_CDNS_7656475930223 $T=20460 5440 0 0 $X=20380 $Y=5190
X200 2 M5_M4_CDNS_7656475930223 $T=22320 4030 0 0 $X=22240 $Y=3780
X201 10 M5_M4_CDNS_7656475930223 $T=24180 3090 0 0 $X=24100 $Y=2840
X202 1 M1_PO_CDNS_7656475930224 $T=930 5440 0 0 $X=830 $Y=5190
X203 3 M1_PO_CDNS_7656475930224 $T=1860 4970 0 0 $X=1760 $Y=4720
X204 2 M1_PO_CDNS_7656475930224 $T=2790 4030 0 0 $X=2690 $Y=3780
X205 6 M1_PO_CDNS_7656475930224 $T=4650 5910 0 0 $X=4550 $Y=5660
X206 1 M1_PO_CDNS_7656475930224 $T=5580 5440 0 0 $X=5480 $Y=5190
X207 3 M1_PO_CDNS_7656475930224 $T=6510 4970 0 0 $X=6410 $Y=4720
X208 2 M1_PO_CDNS_7656475930224 $T=7440 4030 0 0 $X=7340 $Y=3780
X209 7 M1_PO_CDNS_7656475930224 $T=8370 3560 0 0 $X=8270 $Y=3310
X210 9 M1_PO_CDNS_7656475930224 $T=10230 6380 0 0 $X=10130 $Y=6130
X211 6 M1_PO_CDNS_7656475930224 $T=11160 5910 0 0 $X=11060 $Y=5660
X212 1 M1_PO_CDNS_7656475930224 $T=12090 5440 0 0 $X=11990 $Y=5190
X213 3 M1_PO_CDNS_7656475930224 $T=13020 4970 0 0 $X=12920 $Y=4720
X214 2 M1_PO_CDNS_7656475930224 $T=13950 4030 0 0 $X=13850 $Y=3780
X215 7 M1_PO_CDNS_7656475930224 $T=14880 3560 0 0 $X=14780 $Y=3310
X216 10 M1_PO_CDNS_7656475930224 $T=15810 3090 0 0 $X=15710 $Y=2840
X217 12 M1_PO_CDNS_7656475930224 $T=17670 6850 0 0 $X=17570 $Y=6600
X218 9 M1_PO_CDNS_7656475930224 $T=18600 6380 0 0 $X=18500 $Y=6130
X219 6 M1_PO_CDNS_7656475930224 $T=19530 5910 0 0 $X=19430 $Y=5660
X220 1 M1_PO_CDNS_7656475930224 $T=20460 5440 0 0 $X=20360 $Y=5190
X221 3 M1_PO_CDNS_7656475930224 $T=21390 4970 0 0 $X=21290 $Y=4720
X222 2 M1_PO_CDNS_7656475930224 $T=22320 4030 0 0 $X=22220 $Y=3780
X223 7 M1_PO_CDNS_7656475930224 $T=23250 3560 0 0 $X=23150 $Y=3310
X224 10 M1_PO_CDNS_7656475930224 $T=24180 3090 0 0 $X=24080 $Y=2840
X225 14 M1_PO_CDNS_7656475930224 $T=25110 2620 0 0 $X=25010 $Y=2370
X226 1 M2_M1_CDNS_7656475930226 $T=80 5580 0 0 $X=0 $Y=5190
X227 16 M2_M1_CDNS_7656475930226 $T=1540 7840 0 0 $X=1460 $Y=7450
X228 6 M2_M1_CDNS_7656475930226 $T=2130 6050 0 0 $X=2050 $Y=5660
X229 16 M2_M1_CDNS_7656475930226 $T=2470 1570 0 0 $X=2390 $Y=1180
X230 17 M2_M1_CDNS_7656475930226 $T=5260 7840 0 0 $X=5180 $Y=7450
X231 17 M2_M1_CDNS_7656475930226 $T=6450 7840 0 0 $X=6370 $Y=7450
X232 17 M2_M1_CDNS_7656475930226 $T=6860 1570 0 0 $X=6780 $Y=1180
X233 9 M2_M1_CDNS_7656475930226 $T=7710 6520 0 0 $X=7630 $Y=6130
X234 17 M2_M1_CDNS_7656475930226 $T=8050 1570 0 0 $X=7970 $Y=1180
X235 18 M2_M1_CDNS_7656475930226 $T=10840 7840 0 0 $X=10760 $Y=7450
X236 18 M2_M1_CDNS_7656475930226 $T=12030 7840 0 0 $X=11950 $Y=7450
X237 18 M2_M1_CDNS_7656475930226 $T=12960 7840 0 0 $X=12880 $Y=7450
X238 18 M2_M1_CDNS_7656475930226 $T=13370 1570 0 0 $X=13290 $Y=1180
X239 18 M2_M1_CDNS_7656475930226 $T=14300 1570 0 0 $X=14220 $Y=1180
X240 18 M2_M1_CDNS_7656475930226 $T=15490 1570 0 0 $X=15410 $Y=1180
X241 12 M2_M1_CDNS_7656475930226 $T=16080 6990 0 0 $X=16000 $Y=6600
X242 19 M2_M1_CDNS_7656475930226 $T=18280 7840 0 0 $X=18200 $Y=7450
X243 19 M2_M1_CDNS_7656475930226 $T=19470 7840 0 0 $X=19390 $Y=7450
X244 19 M2_M1_CDNS_7656475930226 $T=20400 7840 0 0 $X=20320 $Y=7450
X245 19 M2_M1_CDNS_7656475930226 $T=21330 7840 0 0 $X=21250 $Y=7450
X246 19 M2_M1_CDNS_7656475930226 $T=21740 1570 0 0 $X=21660 $Y=1180
X247 19 M2_M1_CDNS_7656475930226 $T=22670 1570 0 0 $X=22590 $Y=1180
X248 19 M2_M1_CDNS_7656475930226 $T=23600 1570 0 0 $X=23520 $Y=1180
X249 19 M2_M1_CDNS_7656475930226 $T=24790 1570 0 0 $X=24710 $Y=1180
X250 16 M7_M6_CDNS_7656475930227 $T=3580 4500 0 0 $X=3360 $Y=4250
X251 17 M7_M6_CDNS_7656475930227 $T=9160 4500 0 0 $X=8940 $Y=4250
X252 18 M7_M6_CDNS_7656475930227 $T=16600 4500 0 0 $X=16380 $Y=4250
X253 19 M7_M6_CDNS_7656475930227 $T=25900 4500 0 0 $X=25680 $Y=4250
X254 16 M6_M5_CDNS_7656475930228 $T=1540 7840 0 0 $X=1460 $Y=7450
X255 16 M6_M5_CDNS_7656475930228 $T=2470 1570 0 0 $X=2390 $Y=1180
X256 17 M6_M5_CDNS_7656475930228 $T=5260 7840 0 0 $X=5180 $Y=7450
X257 17 M6_M5_CDNS_7656475930228 $T=6450 7840 0 0 $X=6370 $Y=7450
X258 17 M6_M5_CDNS_7656475930228 $T=6860 1570 0 0 $X=6780 $Y=1180
X259 17 M6_M5_CDNS_7656475930228 $T=8050 1570 0 0 $X=7970 $Y=1180
X260 18 M6_M5_CDNS_7656475930228 $T=10840 7840 0 0 $X=10760 $Y=7450
X261 18 M6_M5_CDNS_7656475930228 $T=12030 7840 0 0 $X=11950 $Y=7450
X262 18 M6_M5_CDNS_7656475930228 $T=12960 7840 0 0 $X=12880 $Y=7450
X263 18 M6_M5_CDNS_7656475930228 $T=13370 1570 0 0 $X=13290 $Y=1180
X264 18 M6_M5_CDNS_7656475930228 $T=14300 1570 0 0 $X=14220 $Y=1180
X265 18 M6_M5_CDNS_7656475930228 $T=15490 1570 0 0 $X=15410 $Y=1180
X266 19 M6_M5_CDNS_7656475930228 $T=18280 7840 0 0 $X=18200 $Y=7450
X267 19 M6_M5_CDNS_7656475930228 $T=19470 7840 0 0 $X=19390 $Y=7450
X268 19 M6_M5_CDNS_7656475930228 $T=20400 7840 0 0 $X=20320 $Y=7450
X269 19 M6_M5_CDNS_7656475930228 $T=21330 7840 0 0 $X=21250 $Y=7450
X270 19 M6_M5_CDNS_7656475930228 $T=21740 1570 0 0 $X=21660 $Y=1180
X271 19 M6_M5_CDNS_7656475930228 $T=22670 1570 0 0 $X=22590 $Y=1180
X272 19 M6_M5_CDNS_7656475930228 $T=23600 1570 0 0 $X=23520 $Y=1180
X273 19 M6_M5_CDNS_7656475930228 $T=24790 1570 0 0 $X=24710 $Y=1180
X274 1 M6_M5_CDNS_7656475930229 $T=80 5580 0 0 $X=0 $Y=5190
X275 6 M6_M5_CDNS_7656475930229 $T=2130 6050 0 0 $X=2050 $Y=5660
X276 9 M6_M5_CDNS_7656475930229 $T=7710 6520 0 0 $X=7630 $Y=6130
X277 12 M6_M5_CDNS_7656475930229 $T=16080 6990 0 0 $X=16000 $Y=6600
X278 1 M3_M2_CDNS_7656475930230 $T=80 5580 0 0 $X=0 $Y=5190
X279 16 M3_M2_CDNS_7656475930230 $T=1540 7840 0 0 $X=1460 $Y=7450
X280 6 M3_M2_CDNS_7656475930230 $T=2130 6050 0 0 $X=2050 $Y=5660
X281 16 M3_M2_CDNS_7656475930230 $T=2470 1570 0 0 $X=2390 $Y=1180
X282 17 M3_M2_CDNS_7656475930230 $T=5260 7840 0 0 $X=5180 $Y=7450
X283 17 M3_M2_CDNS_7656475930230 $T=6450 7840 0 0 $X=6370 $Y=7450
X284 17 M3_M2_CDNS_7656475930230 $T=6860 1570 0 0 $X=6780 $Y=1180
X285 9 M3_M2_CDNS_7656475930230 $T=7710 6520 0 0 $X=7630 $Y=6130
X286 17 M3_M2_CDNS_7656475930230 $T=8050 1570 0 0 $X=7970 $Y=1180
X287 18 M3_M2_CDNS_7656475930230 $T=10840 7840 0 0 $X=10760 $Y=7450
X288 18 M3_M2_CDNS_7656475930230 $T=12030 7840 0 0 $X=11950 $Y=7450
X289 18 M3_M2_CDNS_7656475930230 $T=12960 7840 0 0 $X=12880 $Y=7450
X290 18 M3_M2_CDNS_7656475930230 $T=13370 1570 0 0 $X=13290 $Y=1180
X291 18 M3_M2_CDNS_7656475930230 $T=14300 1570 0 0 $X=14220 $Y=1180
X292 18 M3_M2_CDNS_7656475930230 $T=15490 1570 0 0 $X=15410 $Y=1180
X293 12 M3_M2_CDNS_7656475930230 $T=16080 6990 0 0 $X=16000 $Y=6600
X294 19 M3_M2_CDNS_7656475930230 $T=18280 7840 0 0 $X=18200 $Y=7450
X295 19 M3_M2_CDNS_7656475930230 $T=19470 7840 0 0 $X=19390 $Y=7450
X296 19 M3_M2_CDNS_7656475930230 $T=20400 7840 0 0 $X=20320 $Y=7450
X297 19 M3_M2_CDNS_7656475930230 $T=21330 7840 0 0 $X=21250 $Y=7450
X298 19 M3_M2_CDNS_7656475930230 $T=21740 1570 0 0 $X=21660 $Y=1180
X299 19 M3_M2_CDNS_7656475930230 $T=22670 1570 0 0 $X=22590 $Y=1180
X300 19 M3_M2_CDNS_7656475930230 $T=23600 1570 0 0 $X=23520 $Y=1180
X301 19 M3_M2_CDNS_7656475930230 $T=24790 1570 0 0 $X=24710 $Y=1180
X302 1 M5_M4_CDNS_7656475930231 $T=80 5580 0 0 $X=0 $Y=5190
X303 16 M5_M4_CDNS_7656475930231 $T=1540 7840 0 0 $X=1460 $Y=7450
X304 6 M5_M4_CDNS_7656475930231 $T=2130 6050 0 0 $X=2050 $Y=5660
X305 16 M5_M4_CDNS_7656475930231 $T=2470 1570 0 0 $X=2390 $Y=1180
X306 17 M5_M4_CDNS_7656475930231 $T=5260 7840 0 0 $X=5180 $Y=7450
X307 17 M5_M4_CDNS_7656475930231 $T=6450 7840 0 0 $X=6370 $Y=7450
X308 17 M5_M4_CDNS_7656475930231 $T=6860 1570 0 0 $X=6780 $Y=1180
X309 9 M5_M4_CDNS_7656475930231 $T=7710 6520 0 0 $X=7630 $Y=6130
X310 17 M5_M4_CDNS_7656475930231 $T=8050 1570 0 0 $X=7970 $Y=1180
X311 18 M5_M4_CDNS_7656475930231 $T=10840 7840 0 0 $X=10760 $Y=7450
X312 18 M5_M4_CDNS_7656475930231 $T=12030 7840 0 0 $X=11950 $Y=7450
X313 18 M5_M4_CDNS_7656475930231 $T=12960 7840 0 0 $X=12880 $Y=7450
X314 18 M5_M4_CDNS_7656475930231 $T=13370 1570 0 0 $X=13290 $Y=1180
X315 18 M5_M4_CDNS_7656475930231 $T=14300 1570 0 0 $X=14220 $Y=1180
X316 18 M5_M4_CDNS_7656475930231 $T=15490 1570 0 0 $X=15410 $Y=1180
X317 12 M5_M4_CDNS_7656475930231 $T=16080 6990 0 0 $X=16000 $Y=6600
X318 19 M5_M4_CDNS_7656475930231 $T=18280 7840 0 0 $X=18200 $Y=7450
X319 19 M5_M4_CDNS_7656475930231 $T=19470 7840 0 0 $X=19390 $Y=7450
X320 19 M5_M4_CDNS_7656475930231 $T=20400 7840 0 0 $X=20320 $Y=7450
X321 19 M5_M4_CDNS_7656475930231 $T=21330 7840 0 0 $X=21250 $Y=7450
X322 19 M5_M4_CDNS_7656475930231 $T=21740 1570 0 0 $X=21660 $Y=1180
X323 19 M5_M4_CDNS_7656475930231 $T=22670 1570 0 0 $X=22590 $Y=1180
X324 19 M5_M4_CDNS_7656475930231 $T=23600 1570 0 0 $X=23520 $Y=1180
X325 19 M5_M4_CDNS_7656475930231 $T=24790 1570 0 0 $X=24710 $Y=1180
X326 4 4 1 16 5 pmos1v_CDNS_765647593028 $T=1030 8610 1 0 $X=610 $Y=8170
X327 20 4 3 16 5 pmos1v_CDNS_765647593028 $T=2050 8610 0 180 $X=1540 $Y=8170
X328 22 4 1 17 5 pmos1v_CDNS_765647593028 $T=5770 8610 0 180 $X=5260 $Y=8170
X329 4 4 18 13 5 pmos1v_CDNS_765647593028 $T=16840 8610 1 0 $X=16420 $Y=8170
X330 29 4 9 19 5 pmos1v_CDNS_765647593028 $T=18790 8610 0 180 $X=18280 $Y=8170
X331 28 4 3 19 5 pmos1v_CDNS_765647593028 $T=21580 8610 0 180 $X=21070 $Y=8170
X332 29 4 10 26 5 pmos1v_CDNS_765647593028 $T=24370 8610 0 180 $X=23860 $Y=8170
X333 5 5 2 16 nmos1v_CDNS_765647593029 $T=2980 1040 0 180 $X=2470 $Y=240
X334 5 5 16 8 nmos1v_CDNS_765647593029 $T=3820 1040 1 0 $X=3400 $Y=240
X335 31 5 1 37 nmos1v_CDNS_765647593029 $T=5680 1040 1 0 $X=5260 $Y=240
X336 37 5 3 17 nmos1v_CDNS_765647593029 $T=6610 1040 1 0 $X=6190 $Y=240
X337 5 5 9 34 nmos1v_CDNS_765647593029 $T=10330 1040 1 0 $X=9910 $Y=240
X338 34 5 6 32 nmos1v_CDNS_765647593029 $T=11260 1040 1 0 $X=10840 $Y=240
X339 32 5 2 18 nmos1v_CDNS_765647593029 $T=14050 1040 1 0 $X=13630 $Y=240
X340 5 5 12 35 nmos1v_CDNS_765647593029 $T=17770 1040 1 0 $X=17350 $Y=240
X341 36 5 6 38 nmos1v_CDNS_765647593029 $T=19630 1040 1 0 $X=19210 $Y=240
X342 38 5 1 39 nmos1v_CDNS_765647593029 $T=20560 1040 1 0 $X=20140 $Y=240
X343 39 5 3 19 nmos1v_CDNS_765647593029 $T=21490 1040 1 0 $X=21070 $Y=240
X344 38 5 2 19 nmos1v_CDNS_765647593029 $T=22420 1040 1 0 $X=22000 $Y=240
X345 35 5 10 19 nmos1v_CDNS_765647593029 $T=24280 1040 1 0 $X=23860 $Y=240
X346 5 5 14 19 nmos1v_CDNS_765647593029 $T=25300 1040 0 180 $X=24790 $Y=240
M0 4 2 20 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M1 8 16 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M2 17 6 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M3 21 3 17 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M4 22 2 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M5 4 7 22 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M6 11 17 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M7 18 9 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M8 23 6 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M9 24 1 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M10 25 3 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M11 24 2 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M12 23 7 24 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M13 4 10 23 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M14 19 12 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M15 26 6 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M16 27 1 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M17 27 2 28 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M18 26 7 27 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930233                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930233 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930233

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656475930234                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656475930234 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656475930234

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656475930235                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656475930235 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656475930235

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930210                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930210 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930211                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930211 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930211

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930212                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930212 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930212

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930213                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930213 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930213

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930214                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930214 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930214

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930215                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930215 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656475930215

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930216                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930216 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930216

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930217                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930217 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930217

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930218                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930218 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930218

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930219                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930219 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930219

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930220                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930220 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930220

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=16
X0 1 M2_M1_CDNS_7656475930211 $T=2220 -7390 0 90 $X=2090 $Y=-7470
X1 1 M2_M1_CDNS_7656475930211 $T=2220 -4680 0 90 $X=2090 $Y=-4760
X2 7 M2_M1_CDNS_7656475930211 $T=4200 -2840 0 90 $X=4070 $Y=-2920
X3 8 M2_M1_CDNS_7656475930211 $T=4570 -3920 0 90 $X=4440 $Y=-4000
X4 8 M1_PO_CDNS_7656475930214 $T=2340 -4370 0 90 $X=2090 $Y=-4470
X5 8 M1_PO_CDNS_7656475930214 $T=2930 -6480 0 90 $X=2680 $Y=-6580
X6 8 M1_PO_CDNS_7656475930214 $T=2950 -5710 0 90 $X=2700 $Y=-5810
X7 4 M1_PO_CDNS_7656475930214 $T=3490 -4140 0 90 $X=3240 $Y=-4240
X8 4 M1_PO_CDNS_7656475930214 $T=3500 -3460 0 90 $X=3250 $Y=-3560
X9 8 M2_M1_CDNS_7656475930216 $T=2340 -4370 0 90 $X=2090 $Y=-4450
X10 8 M2_M1_CDNS_7656475930216 $T=2930 -6480 0 90 $X=2680 $Y=-6560
X11 8 M2_M1_CDNS_7656475930216 $T=2950 -5710 0 90 $X=2700 $Y=-5790
X12 4 M2_M1_CDNS_7656475930216 $T=3490 -4140 0 90 $X=3240 $Y=-4220
X13 4 M2_M1_CDNS_7656475930216 $T=3500 -3460 0 90 $X=3250 $Y=-3540
X14 9 M2_M1_CDNS_7656475930216 $T=5640 -5920 0 90 $X=5390 $Y=-6000
X15 9 M2_M1_CDNS_7656475930216 $T=5640 -5080 0 90 $X=5390 $Y=-5160
X16 9 M2_M1_CDNS_7656475930216 $T=5640 -4300 0 90 $X=5390 $Y=-4380
X17 6 6 4 8 2 pmos1v_CDNS_765647593020 $T=5520 -3500 0 270 $X=5320 $Y=-4010
X18 6 6 5 7 2 pmos1v_CDNS_765647593020 $T=5520 -2570 0 270 $X=5320 $Y=-3080
X19 2 2 4 8 nmos1v_CDNS_765647593021 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X20 2 2 5 7 nmos1v_CDNS_765647593021 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X21 10 M2_M1_CDNS_7656475930233 $T=1300 -5710 0 90 $X=1170 $Y=-5840
X22 10 M2_M1_CDNS_7656475930233 $T=1300 -4270 0 90 $X=1170 $Y=-4400
X23 4 M2_M1_CDNS_7656475930234 $T=3500 -4810 0 0 $X=3250 $Y=-4940
X24 4 M2_M1_CDNS_7656475930234 $T=3500 -1930 0 0 $X=3250 $Y=-2060
X25 7 M2_M1_CDNS_7656475930234 $T=4210 -6730 0 0 $X=3960 $Y=-6860
X26 7 M2_M1_CDNS_7656475930234 $T=4210 -5370 0 0 $X=3960 $Y=-5500
X27 8 M2_M1_CDNS_7656475930234 $T=4540 -5740 0 0 $X=4290 $Y=-5870
X28 5 M2_M1_CDNS_7656475930234 $T=4960 -4960 0 0 $X=4710 $Y=-5090
X29 5 M2_M1_CDNS_7656475930234 $T=4960 -2500 0 0 $X=4710 $Y=-2630
X30 4 M1_PO_CDNS_7656475930235 $T=3500 -4810 0 0 $X=3260 $Y=-4910
X31 7 M1_PO_CDNS_7656475930235 $T=4210 -6730 0 0 $X=3970 $Y=-6830
X32 7 M1_PO_CDNS_7656475930235 $T=4210 -5370 0 0 $X=3970 $Y=-5470
X33 8 M1_PO_CDNS_7656475930235 $T=4540 -5740 0 0 $X=4300 $Y=-5840
X34 5 M1_PO_CDNS_7656475930235 $T=4960 -4960 0 0 $X=4720 $Y=-5060
X35 5 M1_PO_CDNS_7656475930235 $T=4960 -2500 0 0 $X=4720 $Y=-2600
X36 1 5 9 2 6 pmos1v_CDNS_7656475930210 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 2 7 3 nmos1v_CDNS_7656475930211 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 9 6 7 2 pmos1v_CDNS_7656475930212 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 6 8 11 2 pmos1v_CDNS_7656475930213 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 3 7 11 2 6 pmos1v_CDNS_7656475930214 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X41 2 3 8 2 nmos1v_CDNS_7656475930215 $T=1570 -6390 0 270 $X=1370 $Y=-6840
X42 10 1 8 2 nmos1v_CDNS_7656475930215 $T=1570 -4430 0 270 $X=1370 $Y=-4880
X43 10 7 2 nmos1v_CDNS_7656475930216 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 4 1 12 2 nmos1v_CDNS_7656475930217 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 2 5 12 nmos1v_CDNS_7656475930218 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 9 8 6 2 pmos1v_CDNS_7656475930219 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 9 4 1 2 6 pmos1v_CDNS_7656475930220 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 2 8 3 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 10 8 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M2 6 4 8 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=5520 $Y=-3590 $dt=1
M3 6 5 7 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5520 $Y=-2660 $dt=1
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MAC                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MAC 99 88 84 78 76 72 68 93 89 85
+ 79 77 73 69 64 92 62 97 86 82
+ 80 74 70 66 3 91 87 83 81 75
+ 71 67 65 63 98 57 55 53 51 49
+ 47 60 58 56 54 52 50 48 46 59
+ 61
** N=291 EP=51 FDC=570
X0 1 M3_M2_CDNS_765647593020 $T=150 23850 0 0 $X=70 $Y=23600
X1 2 M3_M2_CDNS_765647593020 $T=5940 23850 0 0 $X=5860 $Y=23600
X2 3 M3_M2_CDNS_765647593020 $T=9840 3330 0 0 $X=9760 $Y=3080
X3 4 M3_M2_CDNS_765647593020 $T=16170 2650 0 0 $X=16090 $Y=2400
X4 5 M3_M2_CDNS_765647593020 $T=16170 23850 0 0 $X=16090 $Y=23600
X5 6 M3_M2_CDNS_765647593020 $T=21750 2650 0 0 $X=21670 $Y=2400
X6 7 M3_M2_CDNS_765647593020 $T=21750 23850 0 0 $X=21670 $Y=23600
X7 8 M3_M2_CDNS_765647593020 $T=26890 2650 0 0 $X=26810 $Y=2400
X8 9 M3_M2_CDNS_765647593020 $T=26890 23850 0 0 $X=26810 $Y=23600
X9 10 M3_M2_CDNS_765647593020 $T=32670 2650 0 0 $X=32590 $Y=2400
X10 11 M3_M2_CDNS_765647593020 $T=32670 23850 0 0 $X=32590 $Y=23600
X11 12 M3_M2_CDNS_765647593020 $T=40090 2650 0 0 $X=40010 $Y=2400
X12 13 M3_M2_CDNS_765647593020 $T=40090 23850 0 0 $X=40010 $Y=23600
X13 14 M3_M2_CDNS_765647593020 $T=48440 2650 0 0 $X=48360 $Y=2400
X14 15 M3_M2_CDNS_765647593020 $T=48440 23850 0 0 $X=48360 $Y=23600
X15 16 M3_M2_CDNS_765647593020 $T=53580 23850 0 0 $X=53500 $Y=23600
X16 1 M4_M3_CDNS_765647593021 $T=150 23850 0 0 $X=70 $Y=23600
X17 2 M4_M3_CDNS_765647593021 $T=5940 23850 0 0 $X=5860 $Y=23600
X18 4 M4_M3_CDNS_765647593021 $T=16170 2650 0 0 $X=16090 $Y=2400
X19 5 M4_M3_CDNS_765647593021 $T=16170 23850 0 0 $X=16090 $Y=23600
X20 6 M4_M3_CDNS_765647593021 $T=21750 2650 0 0 $X=21670 $Y=2400
X21 7 M4_M3_CDNS_765647593021 $T=21750 23850 0 0 $X=21670 $Y=23600
X22 8 M4_M3_CDNS_765647593021 $T=26890 2650 0 0 $X=26810 $Y=2400
X23 9 M4_M3_CDNS_765647593021 $T=26890 23850 0 0 $X=26810 $Y=23600
X24 10 M4_M3_CDNS_765647593021 $T=32670 2650 0 0 $X=32590 $Y=2400
X25 11 M4_M3_CDNS_765647593021 $T=32670 23850 0 0 $X=32590 $Y=23600
X26 12 M4_M3_CDNS_765647593021 $T=40090 2650 0 0 $X=40010 $Y=2400
X27 13 M4_M3_CDNS_765647593021 $T=40090 23850 0 0 $X=40010 $Y=23600
X28 14 M4_M3_CDNS_765647593021 $T=48440 2650 0 0 $X=48360 $Y=2400
X29 15 M4_M3_CDNS_765647593021 $T=48440 23850 0 0 $X=48360 $Y=23600
X30 16 M4_M3_CDNS_765647593021 $T=53580 23850 0 0 $X=53500 $Y=23600
X31 1 M5_M4_CDNS_765647593022 $T=150 23850 0 0 $X=70 $Y=23600
X32 2 M5_M4_CDNS_765647593022 $T=5940 23850 0 0 $X=5860 $Y=23600
X33 4 M5_M4_CDNS_765647593022 $T=16170 2650 0 0 $X=16090 $Y=2400
X34 5 M5_M4_CDNS_765647593022 $T=16170 23850 0 0 $X=16090 $Y=23600
X35 6 M5_M4_CDNS_765647593022 $T=21750 2650 0 0 $X=21670 $Y=2400
X36 7 M5_M4_CDNS_765647593022 $T=21750 23850 0 0 $X=21670 $Y=23600
X37 8 M5_M4_CDNS_765647593022 $T=26890 2650 0 0 $X=26810 $Y=2400
X38 9 M5_M4_CDNS_765647593022 $T=26890 23850 0 0 $X=26810 $Y=23600
X39 10 M5_M4_CDNS_765647593022 $T=32670 2650 0 0 $X=32590 $Y=2400
X40 11 M5_M4_CDNS_765647593022 $T=32670 23850 0 0 $X=32590 $Y=23600
X41 12 M5_M4_CDNS_765647593022 $T=40090 2650 0 0 $X=40010 $Y=2400
X42 13 M5_M4_CDNS_765647593022 $T=40090 23850 0 0 $X=40010 $Y=23600
X43 14 M5_M4_CDNS_765647593022 $T=48440 2650 0 0 $X=48360 $Y=2400
X44 15 M5_M4_CDNS_765647593022 $T=48440 23850 0 0 $X=48360 $Y=23600
X45 16 M5_M4_CDNS_765647593022 $T=53580 23850 0 0 $X=53500 $Y=23600
X46 1 M6_M5_CDNS_765647593023 $T=150 23850 0 0 $X=70 $Y=23600
X47 2 M6_M5_CDNS_765647593023 $T=5940 23850 0 0 $X=5860 $Y=23600
X48 4 M6_M5_CDNS_765647593023 $T=16170 2650 0 0 $X=16090 $Y=2400
X49 5 M6_M5_CDNS_765647593023 $T=16170 23850 0 0 $X=16090 $Y=23600
X50 6 M6_M5_CDNS_765647593023 $T=21750 2650 0 0 $X=21670 $Y=2400
X51 7 M6_M5_CDNS_765647593023 $T=21750 23850 0 0 $X=21670 $Y=23600
X52 8 M6_M5_CDNS_765647593023 $T=26890 2650 0 0 $X=26810 $Y=2400
X53 9 M6_M5_CDNS_765647593023 $T=26890 23850 0 0 $X=26810 $Y=23600
X54 10 M6_M5_CDNS_765647593023 $T=32670 2650 0 0 $X=32590 $Y=2400
X55 11 M6_M5_CDNS_765647593023 $T=32670 23850 0 0 $X=32590 $Y=23600
X56 12 M6_M5_CDNS_765647593023 $T=40090 2650 0 0 $X=40010 $Y=2400
X57 13 M6_M5_CDNS_765647593023 $T=40090 23850 0 0 $X=40010 $Y=23600
X58 14 M6_M5_CDNS_765647593023 $T=48440 2650 0 0 $X=48360 $Y=2400
X59 15 M6_M5_CDNS_765647593023 $T=48440 23850 0 0 $X=48360 $Y=23600
X60 16 M6_M5_CDNS_765647593023 $T=53580 23850 0 0 $X=53500 $Y=23600
X61 17 M3_M2_CDNS_765647593024 $T=560 24410 0 0 $X=480 $Y=24160
X62 18 M3_M2_CDNS_765647593024 $T=9840 24410 0 0 $X=9760 $Y=24160
X63 19 M3_M2_CDNS_765647593024 $T=17280 3210 0 0 $X=17200 $Y=2960
X64 20 M3_M2_CDNS_765647593024 $T=17280 24410 0 0 $X=17200 $Y=24160
X65 21 M3_M2_CDNS_765647593024 $T=22860 3210 0 0 $X=22780 $Y=2960
X66 22 M3_M2_CDNS_765647593024 $T=22860 24410 0 0 $X=22780 $Y=24160
X67 23 M3_M2_CDNS_765647593024 $T=27230 3210 0 0 $X=27150 $Y=2960
X68 24 M3_M2_CDNS_765647593024 $T=27230 24410 0 0 $X=27150 $Y=24160
X69 25 M3_M2_CDNS_765647593024 $T=36530 3210 0 0 $X=36450 $Y=2960
X70 26 M3_M2_CDNS_765647593024 $T=36530 24410 0 0 $X=36450 $Y=24160
X71 27 M3_M2_CDNS_765647593024 $T=43970 3210 0 0 $X=43890 $Y=2960
X72 28 M3_M2_CDNS_765647593024 $T=43970 24410 0 0 $X=43890 $Y=24160
X73 29 M3_M2_CDNS_765647593024 $T=49550 3210 0 0 $X=49470 $Y=2960
X74 30 M3_M2_CDNS_765647593024 $T=49550 24410 0 0 $X=49470 $Y=24160
X75 17 M4_M3_CDNS_765647593025 $T=560 24410 0 0 $X=480 $Y=24160
X76 3 M4_M3_CDNS_765647593025 $T=9840 3330 0 0 $X=9760 $Y=3080
X77 18 M4_M3_CDNS_765647593025 $T=9840 24410 0 0 $X=9760 $Y=24160
X78 19 M4_M3_CDNS_765647593025 $T=17280 3210 0 0 $X=17200 $Y=2960
X79 20 M4_M3_CDNS_765647593025 $T=17280 24410 0 0 $X=17200 $Y=24160
X80 21 M4_M3_CDNS_765647593025 $T=22860 3210 0 0 $X=22780 $Y=2960
X81 22 M4_M3_CDNS_765647593025 $T=22860 24410 0 0 $X=22780 $Y=24160
X82 23 M4_M3_CDNS_765647593025 $T=27230 3210 0 0 $X=27150 $Y=2960
X83 24 M4_M3_CDNS_765647593025 $T=27230 24410 0 0 $X=27150 $Y=24160
X84 25 M4_M3_CDNS_765647593025 $T=36530 3210 0 0 $X=36450 $Y=2960
X85 26 M4_M3_CDNS_765647593025 $T=36530 24410 0 0 $X=36450 $Y=24160
X86 27 M4_M3_CDNS_765647593025 $T=43970 3210 0 0 $X=43890 $Y=2960
X87 28 M4_M3_CDNS_765647593025 $T=43970 24410 0 0 $X=43890 $Y=24160
X88 29 M4_M3_CDNS_765647593025 $T=49550 3210 0 0 $X=49470 $Y=2960
X89 30 M4_M3_CDNS_765647593025 $T=49550 24410 0 0 $X=49470 $Y=24160
X90 31 M3_M2_CDNS_765647593026 $T=9340 41110 0 0 $X=9120 $Y=40860
X91 32 M3_M2_CDNS_765647593026 $T=18130 19910 0 0 $X=17910 $Y=19660
X92 33 M3_M2_CDNS_765647593026 $T=18130 41110 0 0 $X=17910 $Y=40860
X93 34 M3_M2_CDNS_765647593026 $T=23720 19910 0 0 $X=23500 $Y=19660
X94 35 M3_M2_CDNS_765647593026 $T=23720 41110 0 0 $X=23500 $Y=40860
X95 36 M3_M2_CDNS_765647593026 $T=26500 19910 0 0 $X=26280 $Y=19660
X96 37 M3_M2_CDNS_765647593026 $T=26500 41110 0 0 $X=26280 $Y=40860
X97 38 M3_M2_CDNS_765647593026 $T=36030 19910 0 0 $X=35810 $Y=19660
X98 39 M3_M2_CDNS_765647593026 $T=36030 41110 0 0 $X=35810 $Y=40860
X99 40 M3_M2_CDNS_765647593026 $T=44820 19910 0 0 $X=44600 $Y=19660
X100 41 M3_M2_CDNS_765647593026 $T=44820 41110 0 0 $X=44600 $Y=40860
X101 42 M3_M2_CDNS_765647593026 $T=50410 19910 0 0 $X=50190 $Y=19660
X102 43 M3_M2_CDNS_765647593026 $T=50410 41110 0 0 $X=50190 $Y=40860
X103 44 M3_M2_CDNS_765647593026 $T=53190 19910 0 0 $X=52970 $Y=19660
X104 45 M3_M2_CDNS_765647593026 $T=53190 41110 0 0 $X=52970 $Y=40860
X105 31 M4_M3_CDNS_765647593027 $T=9340 41110 0 0 $X=9120 $Y=40860
X106 32 M4_M3_CDNS_765647593027 $T=18130 19910 0 0 $X=17910 $Y=19660
X107 33 M4_M3_CDNS_765647593027 $T=18130 41110 0 0 $X=17910 $Y=40860
X108 34 M4_M3_CDNS_765647593027 $T=23720 19910 0 0 $X=23500 $Y=19660
X109 35 M4_M3_CDNS_765647593027 $T=23720 41110 0 0 $X=23500 $Y=40860
X110 36 M4_M3_CDNS_765647593027 $T=26500 19910 0 0 $X=26280 $Y=19660
X111 37 M4_M3_CDNS_765647593027 $T=26500 41110 0 0 $X=26280 $Y=40860
X112 38 M4_M3_CDNS_765647593027 $T=36030 19910 0 0 $X=35810 $Y=19660
X113 39 M4_M3_CDNS_765647593027 $T=36030 41110 0 0 $X=35810 $Y=40860
X114 40 M4_M3_CDNS_765647593027 $T=44820 19910 0 0 $X=44600 $Y=19660
X115 41 M4_M3_CDNS_765647593027 $T=44820 41110 0 0 $X=44600 $Y=40860
X116 42 M4_M3_CDNS_765647593027 $T=50410 19910 0 0 $X=50190 $Y=19660
X117 43 M4_M3_CDNS_765647593027 $T=50410 41110 0 0 $X=50190 $Y=40860
X118 44 M4_M3_CDNS_765647593027 $T=53190 19910 0 0 $X=52970 $Y=19660
X119 45 M4_M3_CDNS_765647593027 $T=53190 41110 0 0 $X=52970 $Y=40860
X120 31 M5_M4_CDNS_765647593028 $T=9340 41110 0 0 $X=9120 $Y=40860
X121 32 M5_M4_CDNS_765647593028 $T=18130 19910 0 0 $X=17910 $Y=19660
X122 33 M5_M4_CDNS_765647593028 $T=18130 41110 0 0 $X=17910 $Y=40860
X123 34 M5_M4_CDNS_765647593028 $T=23720 19910 0 0 $X=23500 $Y=19660
X124 35 M5_M4_CDNS_765647593028 $T=23720 41110 0 0 $X=23500 $Y=40860
X125 36 M5_M4_CDNS_765647593028 $T=26500 19910 0 0 $X=26280 $Y=19660
X126 37 M5_M4_CDNS_765647593028 $T=26500 41110 0 0 $X=26280 $Y=40860
X127 38 M5_M4_CDNS_765647593028 $T=36030 19910 0 0 $X=35810 $Y=19660
X128 39 M5_M4_CDNS_765647593028 $T=36030 41110 0 0 $X=35810 $Y=40860
X129 40 M5_M4_CDNS_765647593028 $T=44820 19910 0 0 $X=44600 $Y=19660
X130 41 M5_M4_CDNS_765647593028 $T=44820 41110 0 0 $X=44600 $Y=40860
X131 42 M5_M4_CDNS_765647593028 $T=50410 19910 0 0 $X=50190 $Y=19660
X132 43 M5_M4_CDNS_765647593028 $T=50410 41110 0 0 $X=50190 $Y=40860
X133 44 M5_M4_CDNS_765647593028 $T=53190 19910 0 0 $X=52970 $Y=19660
X134 45 M5_M4_CDNS_765647593028 $T=53190 41110 0 0 $X=52970 $Y=40860
X135 31 M6_M5_CDNS_765647593029 $T=9340 41110 0 0 $X=9120 $Y=40860
X136 32 M6_M5_CDNS_765647593029 $T=18130 19910 0 0 $X=17910 $Y=19660
X137 33 M6_M5_CDNS_765647593029 $T=18130 41110 0 0 $X=17910 $Y=40860
X138 34 M6_M5_CDNS_765647593029 $T=23720 19910 0 0 $X=23500 $Y=19660
X139 35 M6_M5_CDNS_765647593029 $T=23720 41110 0 0 $X=23500 $Y=40860
X140 36 M6_M5_CDNS_765647593029 $T=26500 19910 0 0 $X=26280 $Y=19660
X141 37 M6_M5_CDNS_765647593029 $T=26500 41110 0 0 $X=26280 $Y=40860
X142 38 M6_M5_CDNS_765647593029 $T=36030 19910 0 0 $X=35810 $Y=19660
X143 39 M6_M5_CDNS_765647593029 $T=36030 41110 0 0 $X=35810 $Y=40860
X144 40 M6_M5_CDNS_765647593029 $T=44820 19910 0 0 $X=44600 $Y=19660
X145 41 M6_M5_CDNS_765647593029 $T=44820 41110 0 0 $X=44600 $Y=40860
X146 42 M6_M5_CDNS_765647593029 $T=50410 19910 0 0 $X=50190 $Y=19660
X147 43 M6_M5_CDNS_765647593029 $T=50410 41110 0 0 $X=50190 $Y=40860
X148 44 M6_M5_CDNS_765647593029 $T=53190 19910 0 0 $X=52970 $Y=19660
X149 45 M6_M5_CDNS_765647593029 $T=53190 41110 0 0 $X=52970 $Y=40860
X150 31 M2_M1_CDNS_7656475930210 $T=9340 41110 0 0 $X=9120 $Y=40860
X151 32 M2_M1_CDNS_7656475930210 $T=18130 19910 0 0 $X=17910 $Y=19660
X152 33 M2_M1_CDNS_7656475930210 $T=18130 41110 0 0 $X=17910 $Y=40860
X153 34 M2_M1_CDNS_7656475930210 $T=23720 19910 0 0 $X=23500 $Y=19660
X154 35 M2_M1_CDNS_7656475930210 $T=23720 41110 0 0 $X=23500 $Y=40860
X155 36 M2_M1_CDNS_7656475930210 $T=26500 19910 0 0 $X=26280 $Y=19660
X156 37 M2_M1_CDNS_7656475930210 $T=26500 41110 0 0 $X=26280 $Y=40860
X157 38 M2_M1_CDNS_7656475930210 $T=36030 19910 0 0 $X=35810 $Y=19660
X158 39 M2_M1_CDNS_7656475930210 $T=36030 41110 0 0 $X=35810 $Y=40860
X159 40 M2_M1_CDNS_7656475930210 $T=44820 19910 0 0 $X=44600 $Y=19660
X160 41 M2_M1_CDNS_7656475930210 $T=44820 41110 0 0 $X=44600 $Y=40860
X161 42 M2_M1_CDNS_7656475930210 $T=50410 19910 0 0 $X=50190 $Y=19660
X162 43 M2_M1_CDNS_7656475930210 $T=50410 41110 0 0 $X=50190 $Y=40860
X163 44 M2_M1_CDNS_7656475930210 $T=53190 19910 0 0 $X=52970 $Y=19660
X164 45 M2_M1_CDNS_7656475930210 $T=53190 41110 0 0 $X=52970 $Y=40860
X165 46 M2_M1_CDNS_7656475930211 $T=4820 41440 0 0 $X=4740 $Y=41310
X166 47 M2_M1_CDNS_7656475930211 $T=13610 20240 0 0 $X=13530 $Y=20110
X167 48 M2_M1_CDNS_7656475930211 $T=13610 41440 0 0 $X=13530 $Y=41310
X168 49 M2_M1_CDNS_7656475930211 $T=19200 20240 0 0 $X=19120 $Y=20110
X169 50 M2_M1_CDNS_7656475930211 $T=19200 41440 0 0 $X=19120 $Y=41310
X170 51 M2_M1_CDNS_7656475930211 $T=31060 20240 0 0 $X=30980 $Y=20110
X171 52 M2_M1_CDNS_7656475930211 $T=31060 41440 0 0 $X=30980 $Y=41310
X172 53 M2_M1_CDNS_7656475930211 $T=31510 20240 0 0 $X=31430 $Y=20110
X173 54 M2_M1_CDNS_7656475930211 $T=31510 41440 0 0 $X=31430 $Y=41310
X174 55 M2_M1_CDNS_7656475930211 $T=40300 20240 0 0 $X=40220 $Y=20110
X175 56 M2_M1_CDNS_7656475930211 $T=40300 41440 0 0 $X=40220 $Y=41310
X176 57 M2_M1_CDNS_7656475930211 $T=45890 20240 0 0 $X=45810 $Y=20110
X177 58 M2_M1_CDNS_7656475930211 $T=45890 41440 0 0 $X=45810 $Y=41310
X178 59 M2_M1_CDNS_7656475930211 $T=57710 20240 0 0 $X=57630 $Y=20110
X179 60 M2_M1_CDNS_7656475930211 $T=57710 41440 0 0 $X=57630 $Y=41310
X180 3 M2_M1_CDNS_7656475930212 $T=9840 3330 0 0 $X=9760 $Y=3080
X181 17 61 62 63 1 163 100 XOR $T=640 25900 1 0 $X=640 $Y=21200
X182 46 61 62 2 64 164 101 XOR $T=4740 40010 1 0 $X=4740 $Y=35310
X183 18 61 62 65 2 165 102 XOR $T=9740 25900 0 180 $X=6020 $Y=21200
X184 19 61 62 66 4 166 103 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X185 20 61 62 67 5 167 104 XOR $T=17180 25900 0 180 $X=13460 $Y=21200
X186 47 61 62 4 68 168 105 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X187 48 61 62 5 69 169 106 XOR $T=13530 40010 1 0 $X=13530 $Y=35310
X188 21 61 62 70 6 170 107 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X189 22 61 62 71 7 171 108 XOR $T=22760 25900 0 180 $X=19040 $Y=21200
X190 49 61 62 6 72 172 109 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X191 50 61 62 7 73 173 110 XOR $T=19120 40010 1 0 $X=19120 $Y=35310
X192 23 61 62 74 8 174 111 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X193 24 61 62 75 9 175 112 XOR $T=26810 25900 0 180 $X=23090 $Y=21200
X194 51 61 62 8 76 176 113 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X195 52 61 62 9 77 177 114 XOR $T=31140 40010 0 180 $X=27420 $Y=35310
X196 53 61 62 10 78 178 115 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X197 54 61 62 11 79 179 116 XOR $T=31430 40010 1 0 $X=31430 $Y=35310
X198 25 61 62 80 10 180 117 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X199 26 61 62 81 11 181 118 XOR $T=36470 25900 0 180 $X=32750 $Y=21200
X200 27 61 62 82 12 182 119 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X201 28 61 62 83 13 183 120 XOR $T=43890 25900 0 180 $X=40170 $Y=21200
X202 55 61 62 12 84 184 121 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X203 56 61 62 13 85 185 122 XOR $T=40220 40010 1 0 $X=40220 $Y=35310
X204 29 61 62 86 14 186 123 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X205 30 61 62 87 15 187 124 XOR $T=49450 25900 0 180 $X=45730 $Y=21200
X206 57 61 62 14 88 188 125 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X207 58 61 62 15 89 189 126 XOR $T=45810 40010 1 0 $X=45810 $Y=35310
X208 90 61 62 91 16 190 127 XOR $T=49650 25900 1 0 $X=49650 $Y=21200
X209 59 61 62 1 92 191 128 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X210 60 61 62 16 93 192 129 XOR $T=57790 40010 0 180 $X=54070 $Y=35310
X211 64 46 61 62 31 130 193 AND $T=3670 43110 0 0 $X=4740 $Y=40010
X212 68 47 61 62 32 131 194 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X213 69 48 61 62 33 132 195 AND $T=12460 43110 0 0 $X=13530 $Y=40010
X214 72 49 61 62 34 133 196 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X215 73 50 61 62 35 134 197 AND $T=18050 43110 0 0 $X=19120 $Y=40010
X216 76 51 61 62 36 135 198 AND $T=32170 21910 1 180 $X=26920 $Y=18810
X217 77 52 61 62 37 136 199 AND $T=32170 43110 1 180 $X=26920 $Y=40010
X218 78 53 61 62 38 137 200 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X219 79 54 61 62 39 138 201 AND $T=30360 43110 0 0 $X=31430 $Y=40010
X220 84 55 61 62 40 139 202 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X221 85 56 61 62 41 140 203 AND $T=39150 43110 0 0 $X=40220 $Y=40010
X222 88 57 61 62 42 141 204 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X223 89 58 61 62 43 142 205 AND $T=44740 43110 0 0 $X=45810 $Y=40010
X224 92 59 61 62 44 143 206 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X225 93 60 61 62 45 144 207 AND $T=58860 43110 1 180 $X=53610 $Y=40010
X226 8 36 23 61 62 6 34 21 4 32
+ 19 94 3 95 96 145 146 147 148 250
+ 252 251 253 254 255 257 258 259 256 208
+ 209 212 213 211 214 215 210 216 217 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X227 9 37 24 61 62 7 35 22 5 33
+ 20 2 18 31 17 149 150 151 152 260
+ 262 261 263 264 265 267 268 269 266 218
+ 219 222 223 221 224 225 220 226 227 4bit_CLA_logic $T=26970 25900 1 180 $X=320 $Y=25900
X228 1 44 17 61 62 14 42 29 12 40
+ 27 10 25 38 23 153 154 155 156 270
+ 272 271 273 274 275 277 278 279 276 228
+ 229 232 233 231 234 235 230 236 237 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
X229 16 45 90 61 62 15 43 30 13 41
+ 28 11 26 39 24 157 158 159 160 280
+ 282 281 283 284 285 287 288 289 286 238
+ 239 242 243 241 244 245 240 246 247 4bit_CLA_logic $T=53660 25900 1 180 $X=27010 $Y=25900
X230 97 62 90 98 99 61 162 161 290 248
+ 291 249 HAdder $T=62720 27380 1 90 $X=53760 $Y=28180
M0 61 148 96 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M1 61 152 17 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=34270 $dt=1
M2 163 17 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=22000 $dt=1
M3 256 95 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M4 266 31 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=34270 $dt=1
M5 63 1 17 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=22000 $dt=1
M6 163 100 63 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=22000 $dt=1
M7 61 1 100 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=22000 $dt=1
M8 164 46 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=36110 $dt=1
M9 130 46 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=41790 $dt=1
M10 61 64 130 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=41790 $dt=1
M11 2 64 46 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=36110 $dt=1
M12 102 2 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=22000 $dt=1
M13 164 101 2 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=36110 $dt=1
M14 65 102 165 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=22000 $dt=1
M15 61 64 101 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=36110 $dt=1
M16 31 130 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=8230 $Y=41600 $dt=1
M17 18 2 65 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=22000 $dt=1
M18 61 18 165 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=22000 $dt=1
M19 103 4 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M20 104 5 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=115.144 scb=0.0588049 scc=0.0138331 $X=13880 $Y=22000 $dt=1
M21 168 47 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M22 169 48 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=36110 $dt=1
M23 131 47 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.29 scb=0.029437 scc=0.00332952 $X=14390 $Y=20590 $dt=1
M24 132 48 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=41790 $dt=1
M25 61 68 131 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=28.0435 scb=0.0261338 scc=0.00329543 $X=14800 $Y=20590 $dt=1
M26 61 69 132 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=41790 $dt=1
M27 66 103 166 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M28 67 104 167 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.854 scb=0.0354545 scc=0.011187 $X=14810 $Y=22000 $dt=1
M29 4 68 47 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M30 5 69 48 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=36110 $dt=1
M31 19 4 66 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M32 20 5 67 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=15740 $Y=22000 $dt=1
M33 168 105 4 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M34 169 106 5 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=36110 $dt=1
M35 61 19 166 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M36 61 20 167 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=16670 $Y=22000 $dt=1
M37 61 68 105 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M38 61 69 106 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=36110 $dt=1
M39 32 131 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=17020 $Y=20400 $dt=1
M40 33 132 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17020 $Y=41600 $dt=1
M41 107 6 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M42 108 7 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=19460 $Y=22000 $dt=1
M43 172 49 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M44 173 50 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=36110 $dt=1
M45 133 49 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=19980 $Y=20590 $dt=1
M46 134 50 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=41790 $dt=1
M47 70 107 170 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M48 61 72 133 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=20390 $Y=20590 $dt=1
M49 71 108 171 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=20390 $Y=22000 $dt=1
M50 61 73 134 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=41790 $dt=1
M51 6 72 49 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M52 7 73 50 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=36110 $dt=1
M53 21 6 70 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M54 22 7 71 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=21320 $Y=22000 $dt=1
M55 172 109 6 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M56 173 110 7 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=36110 $dt=1
M57 61 21 170 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M58 61 22 171 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=22250 $Y=22000 $dt=1
M59 61 72 109 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M60 61 73 110 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=36110 $dt=1
M61 34 133 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=22610 $Y=20400 $dt=1
M62 35 134 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22610 $Y=41600 $dt=1
M63 111 8 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M64 112 9 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=23510 $Y=22000 $dt=1
M65 74 111 174 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M66 75 112 175 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=24440 $Y=22000 $dt=1
M67 23 8 74 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M68 24 9 75 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=25370 $Y=22000 $dt=1
M69 61 23 174 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M70 61 24 175 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=26300 $Y=22000 $dt=1
M71 61 156 23 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M72 61 160 24 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=34270 $dt=1
M73 61 135 36 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=27520 $Y=20400 $dt=1
M74 61 136 37 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27520 $Y=41600 $dt=1
M75 113 76 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M76 114 77 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=36110 $dt=1
M77 276 38 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M78 286 39 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=34270 $dt=1
M79 8 113 176 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M80 9 114 177 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=36110 $dt=1
M81 51 76 8 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M82 52 77 9 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=36110 $dt=1
M83 135 76 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=29740 $Y=20590 $dt=1
M84 136 77 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29740 $Y=41790 $dt=1
M85 61 51 135 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=30150 $Y=20590 $dt=1
M86 61 52 136 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30150 $Y=41790 $dt=1
M87 61 51 176 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M88 61 52 177 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=36110 $dt=1
M89 178 53 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M90 179 54 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=36110 $dt=1
M91 137 53 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32290 $Y=20590 $dt=1
M92 138 54 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=41790 $dt=1
M93 61 78 137 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32700 $Y=20590 $dt=1
M94 61 79 138 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=41790 $dt=1
M95 10 78 53 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M96 11 79 54 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=36110 $dt=1
M97 117 10 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M98 118 11 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=33170 $Y=22000 $dt=1
M99 178 115 10 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M100 179 116 11 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=36110 $dt=1
M101 80 117 180 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M102 81 118 181 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=34100 $Y=22000 $dt=1
M103 61 78 115 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M104 61 79 116 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=36110 $dt=1
M105 38 137 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=34920 $Y=20400 $dt=1
M106 39 138 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=34920 $Y=41600 $dt=1
M107 25 10 80 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M108 26 11 81 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35030 $Y=22000 $dt=1
M109 61 25 180 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M110 61 26 181 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35960 $Y=22000 $dt=1
M111 119 12 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M112 120 13 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=40590 $Y=22000 $dt=1
M113 184 55 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M114 185 56 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=36110 $dt=1
M115 139 55 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41080 $Y=20590 $dt=1
M116 140 56 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=41790 $dt=1
M117 61 84 139 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41490 $Y=20590 $dt=1
M118 61 85 140 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=41790 $dt=1
M119 82 119 182 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M120 83 120 183 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=41520 $Y=22000 $dt=1
M121 12 84 55 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M122 13 85 56 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=36110 $dt=1
M123 27 12 82 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M124 28 13 83 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=42450 $Y=22000 $dt=1
M125 184 121 12 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M126 185 122 13 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=36110 $dt=1
M127 61 27 182 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M128 61 28 183 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=43380 $Y=22000 $dt=1
M129 61 84 121 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M130 61 85 122 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=36110 $dt=1
M131 40 139 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=43710 $Y=20400 $dt=1
M132 41 140 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=43710 $Y=41600 $dt=1
M133 123 14 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M134 124 15 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=46150 $Y=22000 $dt=1
M135 188 57 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M136 189 58 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=36110 $dt=1
M137 141 57 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=46670 $Y=20590 $dt=1
M138 142 58 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=41790 $dt=1
M139 86 123 186 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M140 61 88 141 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=47080 $Y=20590 $dt=1
M141 87 124 187 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=47080 $Y=22000 $dt=1
M142 61 89 142 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=41790 $dt=1
M143 14 88 57 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M144 15 89 58 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=36110 $dt=1
M145 29 14 86 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=48010 $Y=800 $dt=1
M146 30 15 87 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48010 $Y=22000 $dt=1
M147 188 125 14 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M148 189 126 15 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=36110 $dt=1
M149 61 29 186 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=48940 $Y=800 $dt=1
M150 61 30 187 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48940 $Y=22000 $dt=1
M151 61 88 125 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M152 61 89 126 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=36110 $dt=1
M153 42 141 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=49300 $Y=20400 $dt=1
M154 43 142 61 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=49300 $Y=41600 $dt=1
M155 190 90 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=50070 $Y=22000 $dt=1
M156 91 16 90 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51000 $Y=22000 $dt=1
M157 190 127 91 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51930 $Y=22000 $dt=1
M158 61 16 127 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=52860 $Y=22000 $dt=1
M159 61 143 44 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=54210 $Y=20400 $dt=1
M160 61 144 45 61 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=54210 $Y=41600 $dt=1
M161 128 92 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M162 129 93 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=36110 $dt=1
M163 1 128 191 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M164 16 129 192 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=36110 $dt=1
M165 59 92 1 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M166 60 93 16 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=36110 $dt=1
M167 143 92 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=29.0043 scb=0.0273456 scc=0.00330147 $X=56430 $Y=20590 $dt=1
M168 144 93 61 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=41790 $dt=1
M169 61 59 143 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=33.5338 scb=0.0350848 scc=0.00355838 $X=56840 $Y=20590 $dt=1
M170 61 60 144 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=41790 $dt=1
M171 61 59 191 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M172 61 60 192 61 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=36110 $dt=1
.ends MAC
