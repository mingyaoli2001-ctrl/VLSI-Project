* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 4bit_CLA_logic                               *
* Netlisted  : Sun Dec  7 11:09:58 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765123794261                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765123794261 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765123794261

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765123794262                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765123794262 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765123794262

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic c0 cout1 cout2 cout3 cout4 g1 g2 g3 g4 gnd
+ p1 p2 p3 p4 vdd
** N=39 EP=15 FDC=56
X297 gnd gnd p1 25 nmos1v_CDNS_765123794261 $T=1030 800 0 0 $X=610 $Y=240
X298 25 gnd c0 2 nmos1v_CDNS_765123794261 $T=1960 800 0 0 $X=1540 $Y=240
X299 gnd gnd p2 26 nmos1v_CDNS_765123794261 $T=4750 800 0 0 $X=4330 $Y=240
X300 26 gnd g1 4 nmos1v_CDNS_765123794261 $T=7540 800 0 0 $X=7120 $Y=240
X301 gnd gnd g2 4 nmos1v_CDNS_765123794261 $T=8560 800 1 180 $X=8050 $Y=240
X302 gnd gnd 4 cout2 nmos1v_CDNS_765123794261 $T=9400 800 0 0 $X=8980 $Y=240
X303 27 gnd p1 28 nmos1v_CDNS_765123794261 $T=12190 800 0 0 $X=11770 $Y=240
X304 28 gnd c0 6 nmos1v_CDNS_765123794261 $T=13120 800 0 0 $X=12700 $Y=240
X305 29 gnd g2 6 nmos1v_CDNS_765123794261 $T=14980 800 0 0 $X=14560 $Y=240
X306 gnd gnd g3 6 nmos1v_CDNS_765123794261 $T=16000 800 1 180 $X=15490 $Y=240
X307 gnd gnd 6 cout3 nmos1v_CDNS_765123794261 $T=16840 800 0 0 $X=16420 $Y=240
X308 30 gnd p3 31 nmos1v_CDNS_765123794261 $T=18700 800 0 0 $X=18280 $Y=240
X309 31 gnd g2 8 nmos1v_CDNS_765123794261 $T=23350 800 0 0 $X=22930 $Y=240
X310 gnd gnd 8 cout4 nmos1v_CDNS_765123794261 $T=26140 800 0 0 $X=25720 $Y=240
X311 gnd gnd g1 2 nmos1v_CDNS_765123794262 $T=2980 1040 0 180 $X=2470 $Y=240
X312 gnd gnd 2 cout1 nmos1v_CDNS_765123794262 $T=3820 1040 1 0 $X=3400 $Y=240
X313 26 gnd p1 32 nmos1v_CDNS_765123794262 $T=5680 1040 1 0 $X=5260 $Y=240
X314 32 gnd c0 4 nmos1v_CDNS_765123794262 $T=6610 1040 1 0 $X=6190 $Y=240
X315 gnd gnd p3 29 nmos1v_CDNS_765123794262 $T=10330 1040 1 0 $X=9910 $Y=240
X316 29 gnd p2 27 nmos1v_CDNS_765123794262 $T=11260 1040 1 0 $X=10840 $Y=240
X317 27 gnd g1 6 nmos1v_CDNS_765123794262 $T=14050 1040 1 0 $X=13630 $Y=240
X318 gnd gnd p4 30 nmos1v_CDNS_765123794262 $T=17770 1040 1 0 $X=17350 $Y=240
X319 31 gnd p2 33 nmos1v_CDNS_765123794262 $T=19630 1040 1 0 $X=19210 $Y=240
X320 33 gnd p1 34 nmos1v_CDNS_765123794262 $T=20560 1040 1 0 $X=20140 $Y=240
X321 34 gnd c0 8 nmos1v_CDNS_765123794262 $T=21490 1040 1 0 $X=21070 $Y=240
X322 33 gnd g1 8 nmos1v_CDNS_765123794262 $T=22420 1040 1 0 $X=22000 $Y=240
X323 30 gnd g3 8 nmos1v_CDNS_765123794262 $T=24280 1040 1 0 $X=23860 $Y=240
X324 gnd gnd g4 8 nmos1v_CDNS_765123794262 $T=25300 1040 0 180 $X=24790 $Y=240
M0 2 p1 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1030 $Y=8370 $dt=1
M1 20 c0 2 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1960 $Y=8370 $dt=1
M2 vdd g1 20 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=2890 $Y=8370 $dt=1
M3 cout1 2 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=3820 $Y=8370 $dt=1
M4 4 p2 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=4750 $Y=8370 $dt=1
M5 21 p1 4 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=5680 $Y=8370 $dt=1
M6 35 c0 4 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=6610 $Y=8370 $dt=1
M7 21 g1 35 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=7540 $Y=8370 $dt=1
M8 vdd g2 21 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=8470 $Y=8370 $dt=1
M9 cout2 4 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=9400 $Y=8370 $dt=1
M10 6 p3 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=10330 $Y=8370 $dt=1
M11 36 p2 6 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=11260 $Y=8370 $dt=1
M12 37 p1 6 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=12190 $Y=8370 $dt=1
M13 38 c0 6 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=13120 $Y=8370 $dt=1
M14 37 g1 38 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=14050 $Y=8370 $dt=1
M15 36 g2 37 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=14980 $Y=8370 $dt=1
M16 vdd g3 36 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=15910 $Y=8370 $dt=1
M17 cout3 6 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=16840 $Y=8370 $dt=1
M18 8 p4 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=17770 $Y=8370 $dt=1
M19 22 p3 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=18700 $Y=8370 $dt=1
M20 24 p2 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=19630 $Y=8370 $dt=1
M21 39 p1 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=20560 $Y=8370 $dt=1
M22 23 c0 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21490 $Y=8370 $dt=1
M23 39 g1 23 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22420 $Y=8370 $dt=1
M24 24 g2 39 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23350 $Y=8370 $dt=1
M25 22 g3 24 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24280 $Y=8370 $dt=1
M26 vdd g4 22 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25210 $Y=8370 $dt=1
M27 cout4 8 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26140 $Y=8370 $dt=1
.ends 4bit_CLA_logic
