* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : WallaceProjectMAC                            *
* Netlisted  : Sat Dec 13 20:20:57 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765675251900                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765675251900 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765675251900

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765675251901                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765675251901 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765675251901

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765675251902                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765675251902 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765675251902

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765675251903                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765675251903 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765675251903

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765675251904                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765675251904 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765675251904

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765675251905                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765675251905 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765675251905

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765675251906                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765675251906 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765675251906

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765675251907                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765675251907 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765675251907

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765675251908                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765675251908 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765675251908

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765675251909                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765675251909 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765675251909

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519010                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519010 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519010

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519011                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519011 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519011

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656752519012                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656752519012 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656752519012

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519013                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519013 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519013

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519014                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519014 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519014

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519017                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519017 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519017

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656752519018                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656752519018 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656752519018

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519019                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519019 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519019

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519020                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519020 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519021                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519021 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519023                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519023 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519025                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519025 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519025

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519026                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519026 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519026

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519027                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519027 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519028                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519028 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519028

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519029                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519029 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519029

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519030                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519030 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519030

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519031                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519031 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519031

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519034                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519034 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519034

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519035                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519035 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519035

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519036                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519036 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519036

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519037                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519037 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519037

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519038                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519038 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519038

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519042                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519042 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519042

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519043                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519043 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519043

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519044                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519044 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519044

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656752519045                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656752519045 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656752519045

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656752519047                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656752519047 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656752519047

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656752519049                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656752519049 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656752519049

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519050                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519050 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656752519051                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656752519051 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656752519051

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519052                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519052 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519052

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519053                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519053 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519053

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519054                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519054 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519054

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519056                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519056 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519056

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519058                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519058 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519058

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519059                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519059 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519059

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656752519060                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656752519060 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656752519060

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519061                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519061 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519061

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656752519068                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656752519068 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656752519068

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519069                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519069 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519069

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765675251906                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765675251906 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765675251906

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765675251907                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765675251907 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765675251907

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519071                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519071 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519071

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656752519072                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656752519072 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656752519072

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765675251908                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765675251908 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765675251908

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765675251909                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765675251909 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765675251909

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519010                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519010 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7656752519010

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519011                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519011 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7656752519011

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519012                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519012 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656752519012

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519013                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519013 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656752519013

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519014                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519014 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656752519014

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519015                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519015 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656752519015

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519016                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519016 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656752519016

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519017                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519017 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7656752519017

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519018                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519018 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656752519018

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=8
X0 1 M2_M1_CDNS_7656752519020 $T=2220 -7390 0 90 $X=2090 $Y=-7470
X1 1 M2_M1_CDNS_7656752519020 $T=2220 -4680 0 90 $X=2090 $Y=-4760
X2 7 M2_M1_CDNS_7656752519020 $T=4200 -2840 0 90 $X=4070 $Y=-2920
X3 8 M2_M1_CDNS_7656752519020 $T=4570 -3920 0 90 $X=4440 $Y=-4000
X4 9 M2_M1_CDNS_7656752519025 $T=1300 -5710 0 90 $X=1170 $Y=-5840
X5 9 M2_M1_CDNS_7656752519025 $T=1300 -4270 0 90 $X=1170 $Y=-4400
X6 8 M1_PO_CDNS_7656752519068 $T=2340 -4370 0 90 $X=2090 $Y=-4470
X7 8 M1_PO_CDNS_7656752519068 $T=2930 -6480 0 90 $X=2680 $Y=-6580
X8 8 M1_PO_CDNS_7656752519068 $T=2950 -5710 0 90 $X=2700 $Y=-5810
X9 4 M1_PO_CDNS_7656752519068 $T=3490 -4140 0 90 $X=3240 $Y=-4240
X10 4 M1_PO_CDNS_7656752519068 $T=3500 -3460 0 90 $X=3250 $Y=-3560
X11 8 M2_M1_CDNS_7656752519069 $T=2340 -4370 0 90 $X=2090 $Y=-4450
X12 8 M2_M1_CDNS_7656752519069 $T=2930 -6480 0 90 $X=2680 $Y=-6560
X13 8 M2_M1_CDNS_7656752519069 $T=2950 -5710 0 90 $X=2700 $Y=-5790
X14 4 M2_M1_CDNS_7656752519069 $T=3490 -4140 0 90 $X=3240 $Y=-4220
X15 4 M2_M1_CDNS_7656752519069 $T=3500 -3460 0 90 $X=3250 $Y=-3540
X16 10 M2_M1_CDNS_7656752519069 $T=5640 -5920 0 90 $X=5390 $Y=-6000
X17 10 M2_M1_CDNS_7656752519069 $T=5640 -5080 0 90 $X=5390 $Y=-5160
X18 10 M2_M1_CDNS_7656752519069 $T=5640 -4300 0 90 $X=5390 $Y=-4380
X19 6 6 4 8 2 pmos1v_CDNS_765675251906 $T=5520 -3500 0 270 $X=5320 $Y=-4010
X20 6 6 5 7 2 pmos1v_CDNS_765675251906 $T=5520 -2570 0 270 $X=5320 $Y=-3080
X21 2 2 4 8 nmos1v_CDNS_765675251907 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X22 2 2 5 7 nmos1v_CDNS_765675251907 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X23 4 M2_M1_CDNS_7656752519071 $T=3500 -4810 0 0 $X=3250 $Y=-4940
X24 4 M2_M1_CDNS_7656752519071 $T=3500 -1930 0 0 $X=3250 $Y=-2060
X25 7 M2_M1_CDNS_7656752519071 $T=4210 -6730 0 0 $X=3960 $Y=-6860
X26 7 M2_M1_CDNS_7656752519071 $T=4210 -5370 0 0 $X=3960 $Y=-5500
X27 8 M2_M1_CDNS_7656752519071 $T=4540 -5740 0 0 $X=4290 $Y=-5870
X28 5 M2_M1_CDNS_7656752519071 $T=4960 -4960 0 0 $X=4710 $Y=-5090
X29 5 M2_M1_CDNS_7656752519071 $T=4960 -2500 0 0 $X=4710 $Y=-2630
X30 4 M1_PO_CDNS_7656752519072 $T=3500 -4810 0 0 $X=3260 $Y=-4910
X31 7 M1_PO_CDNS_7656752519072 $T=4210 -6730 0 0 $X=3970 $Y=-6830
X32 7 M1_PO_CDNS_7656752519072 $T=4210 -5370 0 0 $X=3970 $Y=-5470
X33 8 M1_PO_CDNS_7656752519072 $T=4540 -5740 0 0 $X=4300 $Y=-5840
X34 5 M1_PO_CDNS_7656752519072 $T=4960 -4960 0 0 $X=4720 $Y=-5060
X35 5 M1_PO_CDNS_7656752519072 $T=4960 -2500 0 0 $X=4720 $Y=-2600
X36 1 5 10 2 6 pmos1v_CDNS_765675251908 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 2 7 3 nmos1v_CDNS_765675251909 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 10 6 7 2 pmos1v_CDNS_7656752519010 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 6 8 11 2 pmos1v_CDNS_7656752519011 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 3 7 11 2 6 pmos1v_CDNS_7656752519012 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X41 2 3 8 2 nmos1v_CDNS_7656752519013 $T=1570 -6390 0 270 $X=1370 $Y=-6840
X42 9 1 8 2 nmos1v_CDNS_7656752519013 $T=1570 -4430 0 270 $X=1370 $Y=-4880
X43 9 7 2 2 nmos1v_CDNS_7656752519014 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 4 1 12 2 nmos1v_CDNS_7656752519015 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 2 5 12 nmos1v_CDNS_7656752519016 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 10 8 6 2 pmos1v_CDNS_7656752519017 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 10 4 1 2 6 pmos1v_CDNS_7656752519018 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 2 8 3 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 2 7 9 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=6.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-5550 $dt=0
M2 9 8 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M3 2 4 8 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-3590 $dt=0
M4 2 5 7 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1580 $Y=-2660 $dt=0
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656752519062                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656752519062 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656752519062

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519063                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519063 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519063

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519064                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519064 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519064

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519065                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519065 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519065

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519066                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519066 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519066

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656752519067                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656752519067 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656752519067

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765675251900                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765675251900 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_765675251900

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765675251901                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765675251901 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765675251901

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765675251902                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765675251902 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_765675251902

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765675251903                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765675251903 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765675251903

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765675251904                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765675251904 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765675251904

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765675251905                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765675251905 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765675251905

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=0
X0 1 M2_M1_CDNS_7656752519020 $T=1510 -2070 0 0 $X=1430 $Y=-2200
X1 1 M2_M1_CDNS_7656752519020 $T=3010 -2070 0 0 $X=2930 $Y=-2200
X2 5 M3_M2_CDNS_7656752519027 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X3 5 M2_M1_CDNS_7656752519028 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X4 2 M1_PO_CDNS_7656752519067 $T=1870 -1670 0 0 $X=1770 $Y=-1790
X5 1 M1_PO_CDNS_7656752519067 $T=2510 -2070 0 0 $X=2410 $Y=-2190
X6 6 M1_PO_CDNS_7656752519067 $T=4500 -2020 0 0 $X=4400 $Y=-2140
X7 4 5 6 nmos1v_CDNS_765675251900 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X8 3 5 6 4 pmos1v_CDNS_765675251901 $T=4560 -1510 0 0 $X=3880 $Y=-1710
X9 4 1 7 nmos1v_CDNS_765675251902 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X10 3 2 6 4 pmos1v_CDNS_765675251903 $T=1930 -1320 0 0 $X=1250 $Y=-1520
X11 3 6 1 4 pmos1v_CDNS_765675251904 $T=2430 -1320 1 180 $X=1980 $Y=-1520
X12 6 2 7 4 nmos1v_CDNS_765675251905 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X0 6 M2_M1_CDNS_7656752519020 $T=690 3330 0 0 $X=610 $Y=3200
X1 1 M2_M1_CDNS_7656752519020 $T=1190 1490 0 0 $X=1110 $Y=1360
X2 1 M2_M1_CDNS_7656752519020 $T=2520 1490 0 0 $X=2440 $Y=1360
X3 6 M2_M1_CDNS_7656752519020 $T=2550 3330 0 0 $X=2470 $Y=3200
X4 4 M5_M4_CDNS_7656752519062 $T=1850 2810 0 90 $X=1600 $Y=2590
X5 4 M4_M3_CDNS_7656752519063 $T=1850 2810 0 90 $X=1600 $Y=2590
X6 4 M3_M2_CDNS_7656752519064 $T=1850 2810 0 90 $X=1600 $Y=2590
X7 4 M2_M1_CDNS_7656752519065 $T=1850 2810 0 90 $X=1600 $Y=2590
X8 4 M6_M5_CDNS_7656752519066 $T=1850 2810 0 90 $X=1600 $Y=2590
X9 7 M1_PO_CDNS_7656752519067 $T=2470 2570 0 0 $X=2370 $Y=2450
X10 1 M1_PO_CDNS_7656752519068 $T=320 1490 0 0 $X=220 $Y=1240
X11 5 M1_PO_CDNS_7656752519068 $T=1540 2050 0 0 $X=1440 $Y=1800
X12 5 M1_PO_CDNS_7656752519068 $T=3400 2050 0 0 $X=3300 $Y=1800
X13 1 M2_M1_CDNS_7656752519069 $T=320 1490 0 0 $X=240 $Y=1240
X14 5 M2_M1_CDNS_7656752519069 $T=1540 2050 0 0 $X=1460 $Y=1800
X15 5 M2_M1_CDNS_7656752519069 $T=3400 2050 0 0 $X=3320 $Y=1800
X16 3 3 1 6 2 pmos1v_CDNS_765675251906 $T=420 3660 0 0 $X=0 $Y=3460
X17 1 3 5 4 2 pmos1v_CDNS_765675251906 $T=1350 3660 0 0 $X=930 $Y=3460
X18 6 3 7 4 2 pmos1v_CDNS_765675251906 $T=2370 3660 1 180 $X=1860 $Y=3460
X19 3 3 5 7 2 pmos1v_CDNS_765675251906 $T=3300 3660 1 180 $X=2790 $Y=3460
X20 2 2 1 6 nmos1v_CDNS_765675251907 $T=420 800 0 0 $X=0 $Y=240
X21 4 2 5 6 nmos1v_CDNS_765675251907 $T=1440 800 1 180 $X=930 $Y=240
X22 4 2 7 1 nmos1v_CDNS_765675251907 $T=2280 800 0 0 $X=1860 $Y=240
X23 2 2 5 7 nmos1v_CDNS_765675251907 $T=3300 800 1 180 $X=2790 $Y=240
M0 6 1 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=420 $Y=800 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1350 $Y=800 $dt=0
M2 1 7 4 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=2280 $Y=800 $dt=0
M3 2 5 7 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=3210 $Y=800 $dt=0
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656752519073                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656752519073 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656752519073

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656752519074                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656752519074 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656752519074

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656752519075                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656752519075 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656752519075

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519076                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519076 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519076

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656752519077                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656752519077 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656752519077

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519079                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519079 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519079

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656752519080                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656752519080 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656752519080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519081                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519081 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519081

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656752519082                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656752519082 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656752519082

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656752519083                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656752519083 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656752519083

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656752519084                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656752519084 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656752519084

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519019                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519019 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656752519019

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519020                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519020 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656752519020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39
*.DEVICECLIMB
** N=39 EP=39 FDC=54
X0 2 M5_M4_CDNS_765675251908 $T=610 4030 0 0 $X=530 $Y=3780
X1 1 M5_M4_CDNS_765675251908 $T=930 5440 0 0 $X=850 $Y=5190
X2 2 M5_M4_CDNS_765675251908 $T=2790 4030 0 0 $X=2710 $Y=3780
X3 1 M5_M4_CDNS_765675251908 $T=5580 5440 0 0 $X=5500 $Y=5190
X4 2 M5_M4_CDNS_765675251908 $T=7440 4030 0 0 $X=7360 $Y=3780
X5 10 M5_M4_CDNS_765675251908 $T=8700 3090 0 0 $X=8620 $Y=2840
X6 9 M5_M4_CDNS_765675251908 $T=10230 6380 0 0 $X=10150 $Y=6130
X7 1 M5_M4_CDNS_765675251908 $T=12090 5440 0 0 $X=12010 $Y=5190
X8 2 M5_M4_CDNS_765675251908 $T=13950 4030 0 0 $X=13870 $Y=3780
X9 10 M5_M4_CDNS_765675251908 $T=15810 3090 0 0 $X=15730 $Y=2840
X10 9 M5_M4_CDNS_765675251908 $T=18600 6380 0 0 $X=18520 $Y=6130
X11 1 M5_M4_CDNS_765675251908 $T=20460 5440 0 0 $X=20380 $Y=5190
X12 2 M5_M4_CDNS_765675251908 $T=22320 4030 0 0 $X=22240 $Y=3780
X13 10 M5_M4_CDNS_765675251908 $T=24180 3090 0 0 $X=24100 $Y=2840
X14 2 M2_M1_CDNS_765675251909 $T=610 4030 0 0 $X=530 $Y=3780
X15 1 M2_M1_CDNS_765675251909 $T=930 5440 0 0 $X=850 $Y=5190
X16 3 M2_M1_CDNS_765675251909 $T=1860 4970 0 0 $X=1780 $Y=4720
X17 2 M2_M1_CDNS_765675251909 $T=2790 4030 0 0 $X=2710 $Y=3780
X18 7 M2_M1_CDNS_765675251909 $T=3110 3560 0 0 $X=3030 $Y=3310
X19 8 M2_M1_CDNS_765675251909 $T=4110 1490 0 0 $X=4030 $Y=1240
X20 6 M2_M1_CDNS_765675251909 $T=4650 5910 0 0 $X=4570 $Y=5660
X21 1 M2_M1_CDNS_765675251909 $T=5580 5440 0 0 $X=5500 $Y=5190
X22 3 M2_M1_CDNS_765675251909 $T=6510 4970 0 0 $X=6430 $Y=4720
X23 2 M2_M1_CDNS_765675251909 $T=7440 4030 0 0 $X=7360 $Y=3780
X24 7 M2_M1_CDNS_765675251909 $T=8370 3560 0 0 $X=8290 $Y=3310
X25 10 M2_M1_CDNS_765675251909 $T=8700 3090 0 0 $X=8620 $Y=2840
X26 11 M2_M1_CDNS_765675251909 $T=9690 1490 0 0 $X=9610 $Y=1240
X27 9 M2_M1_CDNS_765675251909 $T=10230 6380 0 0 $X=10150 $Y=6130
X28 6 M2_M1_CDNS_765675251909 $T=11160 5910 0 0 $X=11080 $Y=5660
X29 1 M2_M1_CDNS_765675251909 $T=12090 5440 0 0 $X=12010 $Y=5190
X30 3 M2_M1_CDNS_765675251909 $T=13020 4970 0 0 $X=12940 $Y=4720
X31 2 M2_M1_CDNS_765675251909 $T=13950 4030 0 0 $X=13870 $Y=3780
X32 7 M2_M1_CDNS_765675251909 $T=14880 3560 0 0 $X=14800 $Y=3310
X33 10 M2_M1_CDNS_765675251909 $T=15810 3090 0 0 $X=15730 $Y=2840
X34 13 M2_M1_CDNS_765675251909 $T=17130 1490 0 0 $X=17050 $Y=1240
X35 14 M2_M1_CDNS_765675251909 $T=17490 2630 0 0 $X=17410 $Y=2380
X36 12 M2_M1_CDNS_765675251909 $T=17670 6850 0 0 $X=17590 $Y=6600
X37 9 M2_M1_CDNS_765675251909 $T=18600 6380 0 0 $X=18520 $Y=6130
X38 6 M2_M1_CDNS_765675251909 $T=19530 5910 0 0 $X=19450 $Y=5660
X39 1 M2_M1_CDNS_765675251909 $T=20460 5440 0 0 $X=20380 $Y=5190
X40 3 M2_M1_CDNS_765675251909 $T=21390 4970 0 0 $X=21310 $Y=4720
X41 2 M2_M1_CDNS_765675251909 $T=22320 4030 0 0 $X=22240 $Y=3780
X42 7 M2_M1_CDNS_765675251909 $T=23250 3560 0 0 $X=23170 $Y=3310
X43 10 M2_M1_CDNS_765675251909 $T=24180 3090 0 0 $X=24100 $Y=2840
X44 14 M2_M1_CDNS_765675251909 $T=25110 2620 0 0 $X=25030 $Y=2370
X45 15 M2_M1_CDNS_765675251909 $T=26430 1490 0 0 $X=26350 $Y=1240
X46 2 M4_M3_CDNS_7656752519010 $T=610 4030 0 0 $X=530 $Y=3780
X47 1 M4_M3_CDNS_7656752519010 $T=930 5440 0 0 $X=850 $Y=5190
X48 2 M4_M3_CDNS_7656752519010 $T=2790 4030 0 0 $X=2710 $Y=3780
X49 1 M4_M3_CDNS_7656752519010 $T=5580 5440 0 0 $X=5500 $Y=5190
X50 2 M4_M3_CDNS_7656752519010 $T=7440 4030 0 0 $X=7360 $Y=3780
X51 10 M4_M3_CDNS_7656752519010 $T=8700 3090 0 0 $X=8620 $Y=2840
X52 9 M4_M3_CDNS_7656752519010 $T=10230 6380 0 0 $X=10150 $Y=6130
X53 1 M4_M3_CDNS_7656752519010 $T=12090 5440 0 0 $X=12010 $Y=5190
X54 2 M4_M3_CDNS_7656752519010 $T=13950 4030 0 0 $X=13870 $Y=3780
X55 10 M4_M3_CDNS_7656752519010 $T=15810 3090 0 0 $X=15730 $Y=2840
X56 9 M4_M3_CDNS_7656752519010 $T=18600 6380 0 0 $X=18520 $Y=6130
X57 1 M4_M3_CDNS_7656752519010 $T=20460 5440 0 0 $X=20380 $Y=5190
X58 2 M4_M3_CDNS_7656752519010 $T=22320 4030 0 0 $X=22240 $Y=3780
X59 10 M4_M3_CDNS_7656752519010 $T=24180 3090 0 0 $X=24100 $Y=2840
X60 2 M3_M2_CDNS_7656752519011 $T=610 4030 0 0 $X=530 $Y=3780
X61 1 M3_M2_CDNS_7656752519011 $T=930 5440 0 0 $X=850 $Y=5190
X62 2 M3_M2_CDNS_7656752519011 $T=2790 4030 0 0 $X=2710 $Y=3780
X63 7 M3_M2_CDNS_7656752519011 $T=3110 3560 0 0 $X=3030 $Y=3310
X64 8 M3_M2_CDNS_7656752519011 $T=4110 1490 0 0 $X=4030 $Y=1240
X65 1 M3_M2_CDNS_7656752519011 $T=5580 5440 0 0 $X=5500 $Y=5190
X66 2 M3_M2_CDNS_7656752519011 $T=7440 4030 0 0 $X=7360 $Y=3780
X67 10 M3_M2_CDNS_7656752519011 $T=8700 3090 0 0 $X=8620 $Y=2840
X68 11 M3_M2_CDNS_7656752519011 $T=9690 1490 0 0 $X=9610 $Y=1240
X69 9 M3_M2_CDNS_7656752519011 $T=10230 6380 0 0 $X=10150 $Y=6130
X70 1 M3_M2_CDNS_7656752519011 $T=12090 5440 0 0 $X=12010 $Y=5190
X71 2 M3_M2_CDNS_7656752519011 $T=13950 4030 0 0 $X=13870 $Y=3780
X72 10 M3_M2_CDNS_7656752519011 $T=15810 3090 0 0 $X=15730 $Y=2840
X73 13 M3_M2_CDNS_7656752519011 $T=17130 1490 0 0 $X=17050 $Y=1240
X74 14 M3_M2_CDNS_7656752519011 $T=17490 2630 0 0 $X=17410 $Y=2380
X75 9 M3_M2_CDNS_7656752519011 $T=18600 6380 0 0 $X=18520 $Y=6130
X76 1 M3_M2_CDNS_7656752519011 $T=20460 5440 0 0 $X=20380 $Y=5190
X77 2 M3_M2_CDNS_7656752519011 $T=22320 4030 0 0 $X=22240 $Y=3780
X78 10 M3_M2_CDNS_7656752519011 $T=24180 3090 0 0 $X=24100 $Y=2840
X79 15 M3_M2_CDNS_7656752519011 $T=26430 1490 0 0 $X=26350 $Y=1240
X80 3 M3_M2_CDNS_7656752519027 $T=250 4970 0 90 $X=0 $Y=4890
X81 3 M3_M2_CDNS_7656752519027 $T=1860 4970 0 0 $X=1780 $Y=4720
X82 6 M3_M2_CDNS_7656752519027 $T=4650 5910 0 0 $X=4570 $Y=5660
X83 3 M3_M2_CDNS_7656752519027 $T=6510 4970 0 0 $X=6430 $Y=4720
X84 7 M3_M2_CDNS_7656752519027 $T=8370 3560 0 0 $X=8290 $Y=3310
X85 6 M3_M2_CDNS_7656752519027 $T=11160 5910 0 0 $X=11080 $Y=5660
X86 3 M3_M2_CDNS_7656752519027 $T=13020 4970 0 0 $X=12940 $Y=4720
X87 7 M3_M2_CDNS_7656752519027 $T=14880 3560 0 0 $X=14800 $Y=3310
X88 12 M3_M2_CDNS_7656752519027 $T=17670 6850 0 0 $X=17590 $Y=6600
X89 6 M3_M2_CDNS_7656752519027 $T=19530 5910 0 0 $X=19450 $Y=5660
X90 3 M3_M2_CDNS_7656752519027 $T=21390 4970 0 0 $X=21310 $Y=4720
X91 7 M3_M2_CDNS_7656752519027 $T=23250 3560 0 0 $X=23170 $Y=3310
X92 14 M3_M2_CDNS_7656752519027 $T=25110 2620 0 0 $X=25030 $Y=2370
X93 3 M2_M1_CDNS_7656752519028 $T=250 4970 0 90 $X=0 $Y=4890
X94 7 M4_M3_CDNS_7656752519036 $T=3110 3560 0 0 $X=3030 $Y=3310
X95 8 M4_M3_CDNS_7656752519036 $T=4110 1490 0 0 $X=4030 $Y=1240
X96 11 M4_M3_CDNS_7656752519036 $T=9690 1490 0 0 $X=9610 $Y=1240
X97 13 M4_M3_CDNS_7656752519036 $T=17130 1490 0 0 $X=17050 $Y=1240
X98 14 M4_M3_CDNS_7656752519036 $T=17490 2630 0 0 $X=17410 $Y=2380
X99 15 M4_M3_CDNS_7656752519036 $T=26430 1490 0 0 $X=26350 $Y=1240
X100 16 M5_M4_CDNS_7656752519062 $T=3580 4500 0 0 $X=3360 $Y=4250
X101 17 M5_M4_CDNS_7656752519062 $T=9160 4500 0 0 $X=8940 $Y=4250
X102 18 M5_M4_CDNS_7656752519062 $T=16600 4500 0 0 $X=16380 $Y=4250
X103 19 M5_M4_CDNS_7656752519062 $T=25900 4500 0 0 $X=25680 $Y=4250
X104 16 M4_M3_CDNS_7656752519063 $T=3580 4500 0 0 $X=3360 $Y=4250
X105 17 M4_M3_CDNS_7656752519063 $T=9160 4500 0 0 $X=8940 $Y=4250
X106 18 M4_M3_CDNS_7656752519063 $T=16600 4500 0 0 $X=16380 $Y=4250
X107 19 M4_M3_CDNS_7656752519063 $T=25900 4500 0 0 $X=25680 $Y=4250
X108 16 M3_M2_CDNS_7656752519064 $T=3580 4500 0 0 $X=3360 $Y=4250
X109 17 M3_M2_CDNS_7656752519064 $T=9160 4500 0 0 $X=8940 $Y=4250
X110 18 M3_M2_CDNS_7656752519064 $T=16600 4500 0 0 $X=16380 $Y=4250
X111 19 M3_M2_CDNS_7656752519064 $T=25900 4500 0 0 $X=25680 $Y=4250
X112 16 M2_M1_CDNS_7656752519065 $T=3580 4500 0 0 $X=3360 $Y=4250
X113 17 M2_M1_CDNS_7656752519065 $T=9160 4500 0 0 $X=8940 $Y=4250
X114 18 M2_M1_CDNS_7656752519065 $T=16600 4500 0 0 $X=16380 $Y=4250
X115 19 M2_M1_CDNS_7656752519065 $T=25900 4500 0 0 $X=25680 $Y=4250
X116 5 5 2 20 4 pmos1v_CDNS_765675251906 $T=2980 8370 1 180 $X=2470 $Y=8170
X117 5 5 16 8 4 pmos1v_CDNS_765675251906 $T=3820 8370 0 0 $X=3400 $Y=8170
X118 5 5 6 17 4 pmos1v_CDNS_765675251906 $T=4750 8370 0 0 $X=4330 $Y=8170
X119 21 5 3 17 4 pmos1v_CDNS_765675251906 $T=6700 8370 1 180 $X=6190 $Y=8170
X120 22 5 2 21 4 pmos1v_CDNS_765675251906 $T=7630 8370 1 180 $X=7120 $Y=8170
X121 5 5 7 22 4 pmos1v_CDNS_765675251906 $T=8560 8370 1 180 $X=8050 $Y=8170
X122 5 5 17 11 4 pmos1v_CDNS_765675251906 $T=9400 8370 0 0 $X=8980 $Y=8170
X123 5 5 9 18 4 pmos1v_CDNS_765675251906 $T=10330 8370 0 0 $X=9910 $Y=8170
X124 23 5 6 18 4 pmos1v_CDNS_765675251906 $T=11350 8370 1 180 $X=10840 $Y=8170
X125 24 5 1 18 4 pmos1v_CDNS_765675251906 $T=12280 8370 1 180 $X=11770 $Y=8170
X126 25 5 3 18 4 pmos1v_CDNS_765675251906 $T=13210 8370 1 180 $X=12700 $Y=8170
X127 24 5 2 25 4 pmos1v_CDNS_765675251906 $T=14140 8370 1 180 $X=13630 $Y=8170
X128 23 5 7 24 4 pmos1v_CDNS_765675251906 $T=15070 8370 1 180 $X=14560 $Y=8170
X129 5 5 10 23 4 pmos1v_CDNS_765675251906 $T=16000 8370 1 180 $X=15490 $Y=8170
X130 5 5 12 19 4 pmos1v_CDNS_765675251906 $T=17770 8370 0 0 $X=17350 $Y=8170
X131 26 5 6 19 4 pmos1v_CDNS_765675251906 $T=19720 8370 1 180 $X=19210 $Y=8170
X132 27 5 1 19 4 pmos1v_CDNS_765675251906 $T=20650 8370 1 180 $X=20140 $Y=8170
X133 27 5 2 28 4 pmos1v_CDNS_765675251906 $T=22510 8370 1 180 $X=22000 $Y=8170
X134 26 5 7 27 4 pmos1v_CDNS_765675251906 $T=23440 8370 1 180 $X=22930 $Y=8170
X135 5 5 14 29 4 pmos1v_CDNS_765675251906 $T=25300 8370 1 180 $X=24790 $Y=8170
X136 5 5 19 15 4 pmos1v_CDNS_765675251906 $T=26140 8370 0 0 $X=25720 $Y=8170
X137 4 4 1 30 nmos1v_CDNS_765675251907 $T=1030 800 0 0 $X=610 $Y=240
X138 30 4 3 16 nmos1v_CDNS_765675251907 $T=1960 800 0 0 $X=1540 $Y=240
X139 4 4 6 31 nmos1v_CDNS_765675251907 $T=4750 800 0 0 $X=4330 $Y=240
X140 31 4 2 17 nmos1v_CDNS_765675251907 $T=7540 800 0 0 $X=7120 $Y=240
X141 4 4 7 17 nmos1v_CDNS_765675251907 $T=8560 800 1 180 $X=8050 $Y=240
X142 4 4 17 11 nmos1v_CDNS_765675251907 $T=9400 800 0 0 $X=8980 $Y=240
X143 32 4 1 33 nmos1v_CDNS_765675251907 $T=12190 800 0 0 $X=11770 $Y=240
X144 33 4 3 18 nmos1v_CDNS_765675251907 $T=13120 800 0 0 $X=12700 $Y=240
X145 34 4 7 18 nmos1v_CDNS_765675251907 $T=14980 800 0 0 $X=14560 $Y=240
X146 4 4 10 18 nmos1v_CDNS_765675251907 $T=16000 800 1 180 $X=15490 $Y=240
X147 4 4 18 13 nmos1v_CDNS_765675251907 $T=16840 800 0 0 $X=16420 $Y=240
X148 35 4 9 36 nmos1v_CDNS_765675251907 $T=18700 800 0 0 $X=18280 $Y=240
X149 36 4 7 19 nmos1v_CDNS_765675251907 $T=23350 800 0 0 $X=22930 $Y=240
X150 4 4 19 15 nmos1v_CDNS_765675251907 $T=26140 800 0 0 $X=25720 $Y=240
X151 1 M4_M3_CDNS_7656752519073 $T=80 5580 0 0 $X=0 $Y=5190
X152 16 M4_M3_CDNS_7656752519073 $T=1540 7840 0 0 $X=1460 $Y=7450
X153 6 M4_M3_CDNS_7656752519073 $T=2130 6050 0 0 $X=2050 $Y=5660
X154 16 M4_M3_CDNS_7656752519073 $T=2470 1570 0 0 $X=2390 $Y=1180
X155 17 M4_M3_CDNS_7656752519073 $T=5260 7840 0 0 $X=5180 $Y=7450
X156 17 M4_M3_CDNS_7656752519073 $T=6450 7840 0 0 $X=6370 $Y=7450
X157 17 M4_M3_CDNS_7656752519073 $T=6860 1570 0 0 $X=6780 $Y=1180
X158 9 M4_M3_CDNS_7656752519073 $T=7710 6520 0 0 $X=7630 $Y=6130
X159 17 M4_M3_CDNS_7656752519073 $T=8050 1570 0 0 $X=7970 $Y=1180
X160 18 M4_M3_CDNS_7656752519073 $T=10840 7840 0 0 $X=10760 $Y=7450
X161 18 M4_M3_CDNS_7656752519073 $T=12030 7840 0 0 $X=11950 $Y=7450
X162 18 M4_M3_CDNS_7656752519073 $T=12960 7840 0 0 $X=12880 $Y=7450
X163 18 M4_M3_CDNS_7656752519073 $T=13370 1570 0 0 $X=13290 $Y=1180
X164 18 M4_M3_CDNS_7656752519073 $T=14300 1570 0 0 $X=14220 $Y=1180
X165 18 M4_M3_CDNS_7656752519073 $T=15490 1570 0 0 $X=15410 $Y=1180
X166 12 M4_M3_CDNS_7656752519073 $T=16080 6990 0 0 $X=16000 $Y=6600
X167 19 M4_M3_CDNS_7656752519073 $T=18280 7840 0 0 $X=18200 $Y=7450
X168 19 M4_M3_CDNS_7656752519073 $T=19470 7840 0 0 $X=19390 $Y=7450
X169 19 M4_M3_CDNS_7656752519073 $T=20400 7840 0 0 $X=20320 $Y=7450
X170 19 M4_M3_CDNS_7656752519073 $T=21330 7840 0 0 $X=21250 $Y=7450
X171 19 M4_M3_CDNS_7656752519073 $T=21740 1570 0 0 $X=21660 $Y=1180
X172 19 M4_M3_CDNS_7656752519073 $T=22670 1570 0 0 $X=22590 $Y=1180
X173 19 M4_M3_CDNS_7656752519073 $T=23600 1570 0 0 $X=23520 $Y=1180
X174 19 M4_M3_CDNS_7656752519073 $T=24790 1570 0 0 $X=24710 $Y=1180
X175 16 M7_M6_CDNS_7656752519074 $T=1540 7840 0 0 $X=1460 $Y=7450
X176 16 M7_M6_CDNS_7656752519074 $T=2470 1570 0 0 $X=2390 $Y=1180
X177 17 M7_M6_CDNS_7656752519074 $T=5260 7840 0 0 $X=5180 $Y=7450
X178 17 M7_M6_CDNS_7656752519074 $T=6450 7840 0 0 $X=6370 $Y=7450
X179 17 M7_M6_CDNS_7656752519074 $T=6860 1570 0 0 $X=6780 $Y=1180
X180 17 M7_M6_CDNS_7656752519074 $T=8050 1570 0 0 $X=7970 $Y=1180
X181 18 M7_M6_CDNS_7656752519074 $T=10840 7840 0 0 $X=10760 $Y=7450
X182 18 M7_M6_CDNS_7656752519074 $T=12030 7840 0 0 $X=11950 $Y=7450
X183 18 M7_M6_CDNS_7656752519074 $T=12960 7840 0 0 $X=12880 $Y=7450
X184 18 M7_M6_CDNS_7656752519074 $T=13370 1570 0 0 $X=13290 $Y=1180
X185 18 M7_M6_CDNS_7656752519074 $T=14300 1570 0 0 $X=14220 $Y=1180
X186 18 M7_M6_CDNS_7656752519074 $T=15490 1570 0 0 $X=15410 $Y=1180
X187 19 M7_M6_CDNS_7656752519074 $T=18280 7840 0 0 $X=18200 $Y=7450
X188 19 M7_M6_CDNS_7656752519074 $T=19470 7840 0 0 $X=19390 $Y=7450
X189 19 M7_M6_CDNS_7656752519074 $T=20400 7840 0 0 $X=20320 $Y=7450
X190 19 M7_M6_CDNS_7656752519074 $T=21330 7840 0 0 $X=21250 $Y=7450
X191 19 M7_M6_CDNS_7656752519074 $T=21740 1570 0 0 $X=21660 $Y=1180
X192 19 M7_M6_CDNS_7656752519074 $T=22670 1570 0 0 $X=22590 $Y=1180
X193 19 M7_M6_CDNS_7656752519074 $T=23600 1570 0 0 $X=23520 $Y=1180
X194 19 M7_M6_CDNS_7656752519074 $T=24790 1570 0 0 $X=24710 $Y=1180
X195 16 M1_PO_CDNS_7656752519075 $T=3580 4500 0 0 $X=3340 $Y=4250
X196 17 M1_PO_CDNS_7656752519075 $T=9160 4500 0 0 $X=8920 $Y=4250
X197 18 M1_PO_CDNS_7656752519075 $T=16600 4500 0 0 $X=16360 $Y=4250
X198 16 M6_M5_CDNS_7656752519076 $T=3580 4500 0 0 $X=3360 $Y=4250
X199 17 M6_M5_CDNS_7656752519076 $T=9160 4500 0 0 $X=8940 $Y=4250
X200 18 M6_M5_CDNS_7656752519076 $T=16600 4500 0 0 $X=16380 $Y=4250
X201 19 M6_M5_CDNS_7656752519076 $T=25900 4500 0 0 $X=25680 $Y=4250
X202 1 M1_PO_CDNS_7656752519077 $T=930 5440 0 0 $X=830 $Y=5190
X203 3 M1_PO_CDNS_7656752519077 $T=1860 4970 0 0 $X=1760 $Y=4720
X204 2 M1_PO_CDNS_7656752519077 $T=2790 4030 0 0 $X=2690 $Y=3780
X205 6 M1_PO_CDNS_7656752519077 $T=4650 5910 0 0 $X=4550 $Y=5660
X206 1 M1_PO_CDNS_7656752519077 $T=5580 5440 0 0 $X=5480 $Y=5190
X207 3 M1_PO_CDNS_7656752519077 $T=6510 4970 0 0 $X=6410 $Y=4720
X208 2 M1_PO_CDNS_7656752519077 $T=7440 4030 0 0 $X=7340 $Y=3780
X209 7 M1_PO_CDNS_7656752519077 $T=8370 3560 0 0 $X=8270 $Y=3310
X210 9 M1_PO_CDNS_7656752519077 $T=10230 6380 0 0 $X=10130 $Y=6130
X211 6 M1_PO_CDNS_7656752519077 $T=11160 5910 0 0 $X=11060 $Y=5660
X212 1 M1_PO_CDNS_7656752519077 $T=12090 5440 0 0 $X=11990 $Y=5190
X213 3 M1_PO_CDNS_7656752519077 $T=13020 4970 0 0 $X=12920 $Y=4720
X214 2 M1_PO_CDNS_7656752519077 $T=13950 4030 0 0 $X=13850 $Y=3780
X215 7 M1_PO_CDNS_7656752519077 $T=14880 3560 0 0 $X=14780 $Y=3310
X216 10 M1_PO_CDNS_7656752519077 $T=15810 3090 0 0 $X=15710 $Y=2840
X217 12 M1_PO_CDNS_7656752519077 $T=17670 6850 0 0 $X=17570 $Y=6600
X218 9 M1_PO_CDNS_7656752519077 $T=18600 6380 0 0 $X=18500 $Y=6130
X219 6 M1_PO_CDNS_7656752519077 $T=19530 5910 0 0 $X=19430 $Y=5660
X220 1 M1_PO_CDNS_7656752519077 $T=20460 5440 0 0 $X=20360 $Y=5190
X221 3 M1_PO_CDNS_7656752519077 $T=21390 4970 0 0 $X=21290 $Y=4720
X222 2 M1_PO_CDNS_7656752519077 $T=22320 4030 0 0 $X=22220 $Y=3780
X223 7 M1_PO_CDNS_7656752519077 $T=23250 3560 0 0 $X=23150 $Y=3310
X224 10 M1_PO_CDNS_7656752519077 $T=24180 3090 0 0 $X=24080 $Y=2840
X225 14 M1_PO_CDNS_7656752519077 $T=25110 2620 0 0 $X=25010 $Y=2370
X226 1 M2_M1_CDNS_7656752519079 $T=80 5580 0 0 $X=0 $Y=5190
X227 16 M2_M1_CDNS_7656752519079 $T=1540 7840 0 0 $X=1460 $Y=7450
X228 6 M2_M1_CDNS_7656752519079 $T=2130 6050 0 0 $X=2050 $Y=5660
X229 16 M2_M1_CDNS_7656752519079 $T=2470 1570 0 0 $X=2390 $Y=1180
X230 17 M2_M1_CDNS_7656752519079 $T=5260 7840 0 0 $X=5180 $Y=7450
X231 17 M2_M1_CDNS_7656752519079 $T=6450 7840 0 0 $X=6370 $Y=7450
X232 17 M2_M1_CDNS_7656752519079 $T=6860 1570 0 0 $X=6780 $Y=1180
X233 9 M2_M1_CDNS_7656752519079 $T=7710 6520 0 0 $X=7630 $Y=6130
X234 17 M2_M1_CDNS_7656752519079 $T=8050 1570 0 0 $X=7970 $Y=1180
X235 18 M2_M1_CDNS_7656752519079 $T=10840 7840 0 0 $X=10760 $Y=7450
X236 18 M2_M1_CDNS_7656752519079 $T=12030 7840 0 0 $X=11950 $Y=7450
X237 18 M2_M1_CDNS_7656752519079 $T=12960 7840 0 0 $X=12880 $Y=7450
X238 18 M2_M1_CDNS_7656752519079 $T=13370 1570 0 0 $X=13290 $Y=1180
X239 18 M2_M1_CDNS_7656752519079 $T=14300 1570 0 0 $X=14220 $Y=1180
X240 18 M2_M1_CDNS_7656752519079 $T=15490 1570 0 0 $X=15410 $Y=1180
X241 12 M2_M1_CDNS_7656752519079 $T=16080 6990 0 0 $X=16000 $Y=6600
X242 19 M2_M1_CDNS_7656752519079 $T=18280 7840 0 0 $X=18200 $Y=7450
X243 19 M2_M1_CDNS_7656752519079 $T=19470 7840 0 0 $X=19390 $Y=7450
X244 19 M2_M1_CDNS_7656752519079 $T=20400 7840 0 0 $X=20320 $Y=7450
X245 19 M2_M1_CDNS_7656752519079 $T=21330 7840 0 0 $X=21250 $Y=7450
X246 19 M2_M1_CDNS_7656752519079 $T=21740 1570 0 0 $X=21660 $Y=1180
X247 19 M2_M1_CDNS_7656752519079 $T=22670 1570 0 0 $X=22590 $Y=1180
X248 19 M2_M1_CDNS_7656752519079 $T=23600 1570 0 0 $X=23520 $Y=1180
X249 19 M2_M1_CDNS_7656752519079 $T=24790 1570 0 0 $X=24710 $Y=1180
X250 16 M7_M6_CDNS_7656752519080 $T=3580 4500 0 0 $X=3360 $Y=4250
X251 17 M7_M6_CDNS_7656752519080 $T=9160 4500 0 0 $X=8940 $Y=4250
X252 18 M7_M6_CDNS_7656752519080 $T=16600 4500 0 0 $X=16380 $Y=4250
X253 19 M7_M6_CDNS_7656752519080 $T=25900 4500 0 0 $X=25680 $Y=4250
X254 16 M6_M5_CDNS_7656752519081 $T=1540 7840 0 0 $X=1460 $Y=7450
X255 16 M6_M5_CDNS_7656752519081 $T=2470 1570 0 0 $X=2390 $Y=1180
X256 17 M6_M5_CDNS_7656752519081 $T=5260 7840 0 0 $X=5180 $Y=7450
X257 17 M6_M5_CDNS_7656752519081 $T=6450 7840 0 0 $X=6370 $Y=7450
X258 17 M6_M5_CDNS_7656752519081 $T=6860 1570 0 0 $X=6780 $Y=1180
X259 17 M6_M5_CDNS_7656752519081 $T=8050 1570 0 0 $X=7970 $Y=1180
X260 18 M6_M5_CDNS_7656752519081 $T=10840 7840 0 0 $X=10760 $Y=7450
X261 18 M6_M5_CDNS_7656752519081 $T=12030 7840 0 0 $X=11950 $Y=7450
X262 18 M6_M5_CDNS_7656752519081 $T=12960 7840 0 0 $X=12880 $Y=7450
X263 18 M6_M5_CDNS_7656752519081 $T=13370 1570 0 0 $X=13290 $Y=1180
X264 18 M6_M5_CDNS_7656752519081 $T=14300 1570 0 0 $X=14220 $Y=1180
X265 18 M6_M5_CDNS_7656752519081 $T=15490 1570 0 0 $X=15410 $Y=1180
X266 19 M6_M5_CDNS_7656752519081 $T=18280 7840 0 0 $X=18200 $Y=7450
X267 19 M6_M5_CDNS_7656752519081 $T=19470 7840 0 0 $X=19390 $Y=7450
X268 19 M6_M5_CDNS_7656752519081 $T=20400 7840 0 0 $X=20320 $Y=7450
X269 19 M6_M5_CDNS_7656752519081 $T=21330 7840 0 0 $X=21250 $Y=7450
X270 19 M6_M5_CDNS_7656752519081 $T=21740 1570 0 0 $X=21660 $Y=1180
X271 19 M6_M5_CDNS_7656752519081 $T=22670 1570 0 0 $X=22590 $Y=1180
X272 19 M6_M5_CDNS_7656752519081 $T=23600 1570 0 0 $X=23520 $Y=1180
X273 19 M6_M5_CDNS_7656752519081 $T=24790 1570 0 0 $X=24710 $Y=1180
X274 1 M6_M5_CDNS_7656752519082 $T=80 5580 0 0 $X=0 $Y=5190
X275 6 M6_M5_CDNS_7656752519082 $T=2130 6050 0 0 $X=2050 $Y=5660
X276 9 M6_M5_CDNS_7656752519082 $T=7710 6520 0 0 $X=7630 $Y=6130
X277 12 M6_M5_CDNS_7656752519082 $T=16080 6990 0 0 $X=16000 $Y=6600
X278 1 M3_M2_CDNS_7656752519083 $T=80 5580 0 0 $X=0 $Y=5190
X279 16 M3_M2_CDNS_7656752519083 $T=1540 7840 0 0 $X=1460 $Y=7450
X280 6 M3_M2_CDNS_7656752519083 $T=2130 6050 0 0 $X=2050 $Y=5660
X281 16 M3_M2_CDNS_7656752519083 $T=2470 1570 0 0 $X=2390 $Y=1180
X282 17 M3_M2_CDNS_7656752519083 $T=5260 7840 0 0 $X=5180 $Y=7450
X283 17 M3_M2_CDNS_7656752519083 $T=6450 7840 0 0 $X=6370 $Y=7450
X284 17 M3_M2_CDNS_7656752519083 $T=6860 1570 0 0 $X=6780 $Y=1180
X285 9 M3_M2_CDNS_7656752519083 $T=7710 6520 0 0 $X=7630 $Y=6130
X286 17 M3_M2_CDNS_7656752519083 $T=8050 1570 0 0 $X=7970 $Y=1180
X287 18 M3_M2_CDNS_7656752519083 $T=10840 7840 0 0 $X=10760 $Y=7450
X288 18 M3_M2_CDNS_7656752519083 $T=12030 7840 0 0 $X=11950 $Y=7450
X289 18 M3_M2_CDNS_7656752519083 $T=12960 7840 0 0 $X=12880 $Y=7450
X290 18 M3_M2_CDNS_7656752519083 $T=13370 1570 0 0 $X=13290 $Y=1180
X291 18 M3_M2_CDNS_7656752519083 $T=14300 1570 0 0 $X=14220 $Y=1180
X292 18 M3_M2_CDNS_7656752519083 $T=15490 1570 0 0 $X=15410 $Y=1180
X293 12 M3_M2_CDNS_7656752519083 $T=16080 6990 0 0 $X=16000 $Y=6600
X294 19 M3_M2_CDNS_7656752519083 $T=18280 7840 0 0 $X=18200 $Y=7450
X295 19 M3_M2_CDNS_7656752519083 $T=19470 7840 0 0 $X=19390 $Y=7450
X296 19 M3_M2_CDNS_7656752519083 $T=20400 7840 0 0 $X=20320 $Y=7450
X297 19 M3_M2_CDNS_7656752519083 $T=21330 7840 0 0 $X=21250 $Y=7450
X298 19 M3_M2_CDNS_7656752519083 $T=21740 1570 0 0 $X=21660 $Y=1180
X299 19 M3_M2_CDNS_7656752519083 $T=22670 1570 0 0 $X=22590 $Y=1180
X300 19 M3_M2_CDNS_7656752519083 $T=23600 1570 0 0 $X=23520 $Y=1180
X301 19 M3_M2_CDNS_7656752519083 $T=24790 1570 0 0 $X=24710 $Y=1180
X302 1 M5_M4_CDNS_7656752519084 $T=80 5580 0 0 $X=0 $Y=5190
X303 16 M5_M4_CDNS_7656752519084 $T=1540 7840 0 0 $X=1460 $Y=7450
X304 6 M5_M4_CDNS_7656752519084 $T=2130 6050 0 0 $X=2050 $Y=5660
X305 16 M5_M4_CDNS_7656752519084 $T=2470 1570 0 0 $X=2390 $Y=1180
X306 17 M5_M4_CDNS_7656752519084 $T=5260 7840 0 0 $X=5180 $Y=7450
X307 17 M5_M4_CDNS_7656752519084 $T=6450 7840 0 0 $X=6370 $Y=7450
X308 17 M5_M4_CDNS_7656752519084 $T=6860 1570 0 0 $X=6780 $Y=1180
X309 9 M5_M4_CDNS_7656752519084 $T=7710 6520 0 0 $X=7630 $Y=6130
X310 17 M5_M4_CDNS_7656752519084 $T=8050 1570 0 0 $X=7970 $Y=1180
X311 18 M5_M4_CDNS_7656752519084 $T=10840 7840 0 0 $X=10760 $Y=7450
X312 18 M5_M4_CDNS_7656752519084 $T=12030 7840 0 0 $X=11950 $Y=7450
X313 18 M5_M4_CDNS_7656752519084 $T=12960 7840 0 0 $X=12880 $Y=7450
X314 18 M5_M4_CDNS_7656752519084 $T=13370 1570 0 0 $X=13290 $Y=1180
X315 18 M5_M4_CDNS_7656752519084 $T=14300 1570 0 0 $X=14220 $Y=1180
X316 18 M5_M4_CDNS_7656752519084 $T=15490 1570 0 0 $X=15410 $Y=1180
X317 12 M5_M4_CDNS_7656752519084 $T=16080 6990 0 0 $X=16000 $Y=6600
X318 19 M5_M4_CDNS_7656752519084 $T=18280 7840 0 0 $X=18200 $Y=7450
X319 19 M5_M4_CDNS_7656752519084 $T=19470 7840 0 0 $X=19390 $Y=7450
X320 19 M5_M4_CDNS_7656752519084 $T=20400 7840 0 0 $X=20320 $Y=7450
X321 19 M5_M4_CDNS_7656752519084 $T=21330 7840 0 0 $X=21250 $Y=7450
X322 19 M5_M4_CDNS_7656752519084 $T=21740 1570 0 0 $X=21660 $Y=1180
X323 19 M5_M4_CDNS_7656752519084 $T=22670 1570 0 0 $X=22590 $Y=1180
X324 19 M5_M4_CDNS_7656752519084 $T=23600 1570 0 0 $X=23520 $Y=1180
X325 19 M5_M4_CDNS_7656752519084 $T=24790 1570 0 0 $X=24710 $Y=1180
X326 5 5 1 16 4 pmos1v_CDNS_7656752519019 $T=1030 8610 1 0 $X=610 $Y=8170
X327 20 5 3 16 4 pmos1v_CDNS_7656752519019 $T=2050 8610 0 180 $X=1540 $Y=8170
X328 22 5 1 17 4 pmos1v_CDNS_7656752519019 $T=5770 8610 0 180 $X=5260 $Y=8170
X329 5 5 18 13 4 pmos1v_CDNS_7656752519019 $T=16840 8610 1 0 $X=16420 $Y=8170
X330 29 5 9 19 4 pmos1v_CDNS_7656752519019 $T=18790 8610 0 180 $X=18280 $Y=8170
X331 28 5 3 19 4 pmos1v_CDNS_7656752519019 $T=21580 8610 0 180 $X=21070 $Y=8170
X332 29 5 10 26 4 pmos1v_CDNS_7656752519019 $T=24370 8610 0 180 $X=23860 $Y=8170
X333 4 4 2 16 nmos1v_CDNS_7656752519020 $T=2980 1040 0 180 $X=2470 $Y=240
X334 4 4 16 8 nmos1v_CDNS_7656752519020 $T=3820 1040 1 0 $X=3400 $Y=240
X335 31 4 1 37 nmos1v_CDNS_7656752519020 $T=5680 1040 1 0 $X=5260 $Y=240
X336 37 4 3 17 nmos1v_CDNS_7656752519020 $T=6610 1040 1 0 $X=6190 $Y=240
X337 4 4 9 34 nmos1v_CDNS_7656752519020 $T=10330 1040 1 0 $X=9910 $Y=240
X338 34 4 6 32 nmos1v_CDNS_7656752519020 $T=11260 1040 1 0 $X=10840 $Y=240
X339 32 4 2 18 nmos1v_CDNS_7656752519020 $T=14050 1040 1 0 $X=13630 $Y=240
X340 4 4 12 35 nmos1v_CDNS_7656752519020 $T=17770 1040 1 0 $X=17350 $Y=240
X341 36 4 6 38 nmos1v_CDNS_7656752519020 $T=19630 1040 1 0 $X=19210 $Y=240
X342 38 4 1 39 nmos1v_CDNS_7656752519020 $T=20560 1040 1 0 $X=20140 $Y=240
X343 39 4 3 19 nmos1v_CDNS_7656752519020 $T=21490 1040 1 0 $X=21070 $Y=240
X344 38 4 2 19 nmos1v_CDNS_7656752519020 $T=22420 1040 1 0 $X=22000 $Y=240
X345 35 4 10 19 nmos1v_CDNS_7656752519020 $T=24280 1040 1 0 $X=23860 $Y=240
X346 4 4 14 19 nmos1v_CDNS_7656752519020 $T=25300 1040 0 180 $X=24790 $Y=240
M0 30 1 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1030 $Y=800 $dt=0
M1 16 3 30 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1960 $Y=800 $dt=0
M2 31 6 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=4750 $Y=800 $dt=0
M3 17 2 31 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=7540 $Y=800 $dt=0
M4 4 7 17 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=8470 $Y=800 $dt=0
M5 11 17 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=9400 $Y=800 $dt=0
M6 33 1 32 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12190 $Y=800 $dt=0
M7 18 3 33 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=13120 $Y=800 $dt=0
M8 18 7 34 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=14980 $Y=800 $dt=0
M9 4 10 18 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=15910 $Y=800 $dt=0
M10 13 18 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=16840 $Y=800 $dt=0
M11 36 9 35 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=18700 $Y=800 $dt=0
M12 19 7 36 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=23350 $Y=800 $dt=0
M13 15 19 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=26140 $Y=800 $dt=0
M14 16 1 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=1030 $Y=8370 $dt=1
M15 20 3 16 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=1960 $Y=8370 $dt=1
M16 5 2 20 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M17 8 16 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M18 17 6 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M19 22 1 17 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=5680 $Y=8370 $dt=1
M20 21 3 17 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M21 22 2 21 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M22 5 7 22 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M23 11 17 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M24 18 9 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M25 23 6 18 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M26 24 1 18 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M27 25 3 18 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M28 24 2 25 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M29 23 7 24 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M30 5 10 23 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M31 13 18 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=16840 $Y=8370 $dt=1
M32 19 12 5 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M33 29 9 19 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=18700 $Y=8370 $dt=1
M34 26 6 19 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M35 27 1 19 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M36 28 3 19 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=21490 $Y=8370 $dt=1
M37 27 2 28 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M38 26 7 27 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
M39 29 10 26 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=24280 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceFinalAdder                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceFinalAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58
** N=164 EP=58 FDC=320
X0 33 M4_M3_CDNS_7656752519010 $T=150 2650 0 0 $X=70 $Y=2400
X1 34 M4_M3_CDNS_7656752519010 $T=5940 2650 0 0 $X=5860 $Y=2400
X2 35 M4_M3_CDNS_7656752519010 $T=16170 2650 0 0 $X=16090 $Y=2400
X3 36 M4_M3_CDNS_7656752519010 $T=21750 2650 0 0 $X=21670 $Y=2400
X4 37 M4_M3_CDNS_7656752519010 $T=26890 2650 0 0 $X=26810 $Y=2400
X5 38 M4_M3_CDNS_7656752519010 $T=32670 2650 0 0 $X=32590 $Y=2400
X6 39 M4_M3_CDNS_7656752519010 $T=40090 2650 0 0 $X=40010 $Y=2400
X7 40 M4_M3_CDNS_7656752519010 $T=48440 2650 0 0 $X=48360 $Y=2400
X8 41 M4_M3_CDNS_7656752519010 $T=53580 2650 0 0 $X=53500 $Y=2400
X9 33 M3_M2_CDNS_7656752519011 $T=150 2650 0 0 $X=70 $Y=2400
X10 34 M3_M2_CDNS_7656752519011 $T=5940 2650 0 0 $X=5860 $Y=2400
X11 35 M3_M2_CDNS_7656752519011 $T=16170 2650 0 0 $X=16090 $Y=2400
X12 36 M3_M2_CDNS_7656752519011 $T=21750 2650 0 0 $X=21670 $Y=2400
X13 37 M3_M2_CDNS_7656752519011 $T=26890 2650 0 0 $X=26810 $Y=2400
X14 38 M3_M2_CDNS_7656752519011 $T=32670 2650 0 0 $X=32590 $Y=2400
X15 39 M3_M2_CDNS_7656752519011 $T=40090 2650 0 0 $X=40010 $Y=2400
X16 40 M3_M2_CDNS_7656752519011 $T=48440 2650 0 0 $X=48360 $Y=2400
X17 41 M3_M2_CDNS_7656752519011 $T=53580 2650 0 0 $X=53500 $Y=2400
X18 2 M2_M1_CDNS_7656752519020 $T=4820 20240 0 0 $X=4740 $Y=20110
X19 9 M2_M1_CDNS_7656752519020 $T=13610 20240 0 0 $X=13530 $Y=20110
X20 11 M2_M1_CDNS_7656752519020 $T=19200 20240 0 0 $X=19120 $Y=20110
X21 16 M2_M1_CDNS_7656752519020 $T=31060 20240 0 0 $X=30980 $Y=20110
X22 18 M2_M1_CDNS_7656752519020 $T=31510 20240 0 0 $X=31430 $Y=20110
X23 22 M2_M1_CDNS_7656752519020 $T=40300 20240 0 0 $X=40220 $Y=20110
X24 25 M2_M1_CDNS_7656752519020 $T=45890 20240 0 0 $X=45810 $Y=20110
X25 28 M2_M1_CDNS_7656752519020 $T=57710 20240 0 0 $X=57630 $Y=20110
X26 42 M3_M2_CDNS_7656752519035 $T=560 3210 0 0 $X=480 $Y=2960
X27 43 M3_M2_CDNS_7656752519035 $T=9840 3210 0 0 $X=9760 $Y=2960
X28 44 M3_M2_CDNS_7656752519035 $T=17280 3210 0 0 $X=17200 $Y=2960
X29 45 M3_M2_CDNS_7656752519035 $T=22860 3210 0 0 $X=22780 $Y=2960
X30 46 M3_M2_CDNS_7656752519035 $T=27230 3210 0 0 $X=27150 $Y=2960
X31 47 M3_M2_CDNS_7656752519035 $T=36530 3210 0 0 $X=36450 $Y=2960
X32 48 M3_M2_CDNS_7656752519035 $T=43970 3210 0 0 $X=43890 $Y=2960
X33 49 M3_M2_CDNS_7656752519035 $T=49550 3210 0 0 $X=49470 $Y=2960
X34 42 M4_M3_CDNS_7656752519036 $T=560 3210 0 0 $X=480 $Y=2960
X35 43 M4_M3_CDNS_7656752519036 $T=9840 3210 0 0 $X=9760 $Y=2960
X36 44 M4_M3_CDNS_7656752519036 $T=17280 3210 0 0 $X=17200 $Y=2960
X37 45 M4_M3_CDNS_7656752519036 $T=22860 3210 0 0 $X=22780 $Y=2960
X38 46 M4_M3_CDNS_7656752519036 $T=27230 3210 0 0 $X=27150 $Y=2960
X39 47 M4_M3_CDNS_7656752519036 $T=36530 3210 0 0 $X=36450 $Y=2960
X40 48 M4_M3_CDNS_7656752519036 $T=43970 3210 0 0 $X=43890 $Y=2960
X41 49 M4_M3_CDNS_7656752519036 $T=49550 3210 0 0 $X=49470 $Y=2960
X42 33 M5_M4_CDNS_7656752519045 $T=150 2650 0 0 $X=70 $Y=2400
X43 34 M5_M4_CDNS_7656752519045 $T=5940 2650 0 0 $X=5860 $Y=2400
X44 35 M5_M4_CDNS_7656752519045 $T=16170 2650 0 0 $X=16090 $Y=2400
X45 36 M5_M4_CDNS_7656752519045 $T=21750 2650 0 0 $X=21670 $Y=2400
X46 37 M5_M4_CDNS_7656752519045 $T=26890 2650 0 0 $X=26810 $Y=2400
X47 38 M5_M4_CDNS_7656752519045 $T=32670 2650 0 0 $X=32590 $Y=2400
X48 39 M5_M4_CDNS_7656752519045 $T=40090 2650 0 0 $X=40010 $Y=2400
X49 40 M5_M4_CDNS_7656752519045 $T=48440 2650 0 0 $X=48360 $Y=2400
X50 41 M5_M4_CDNS_7656752519045 $T=53580 2650 0 0 $X=53500 $Y=2400
X51 33 M6_M5_CDNS_7656752519053 $T=150 2650 0 0 $X=70 $Y=2400
X52 34 M6_M5_CDNS_7656752519053 $T=5940 2650 0 0 $X=5860 $Y=2400
X53 35 M6_M5_CDNS_7656752519053 $T=16170 2650 0 0 $X=16090 $Y=2400
X54 36 M6_M5_CDNS_7656752519053 $T=21750 2650 0 0 $X=21670 $Y=2400
X55 37 M6_M5_CDNS_7656752519053 $T=26890 2650 0 0 $X=26810 $Y=2400
X56 38 M6_M5_CDNS_7656752519053 $T=32670 2650 0 0 $X=32590 $Y=2400
X57 39 M6_M5_CDNS_7656752519053 $T=40090 2650 0 0 $X=40010 $Y=2400
X58 40 M6_M5_CDNS_7656752519053 $T=48440 2650 0 0 $X=48360 $Y=2400
X59 41 M6_M5_CDNS_7656752519053 $T=53580 2650 0 0 $X=53500 $Y=2400
X60 50 M5_M4_CDNS_7656752519062 $T=9340 19910 0 0 $X=9120 $Y=19660
X61 51 M5_M4_CDNS_7656752519062 $T=18130 19910 0 0 $X=17910 $Y=19660
X62 52 M5_M4_CDNS_7656752519062 $T=23720 19910 0 0 $X=23500 $Y=19660
X63 53 M5_M4_CDNS_7656752519062 $T=26500 19910 0 0 $X=26280 $Y=19660
X64 54 M5_M4_CDNS_7656752519062 $T=36030 19910 0 0 $X=35810 $Y=19660
X65 55 M5_M4_CDNS_7656752519062 $T=44820 19910 0 0 $X=44600 $Y=19660
X66 56 M5_M4_CDNS_7656752519062 $T=50410 19910 0 0 $X=50190 $Y=19660
X67 57 M5_M4_CDNS_7656752519062 $T=53190 19910 0 0 $X=52970 $Y=19660
X68 50 M4_M3_CDNS_7656752519063 $T=9340 19910 0 0 $X=9120 $Y=19660
X69 51 M4_M3_CDNS_7656752519063 $T=18130 19910 0 0 $X=17910 $Y=19660
X70 52 M4_M3_CDNS_7656752519063 $T=23720 19910 0 0 $X=23500 $Y=19660
X71 53 M4_M3_CDNS_7656752519063 $T=26500 19910 0 0 $X=26280 $Y=19660
X72 54 M4_M3_CDNS_7656752519063 $T=36030 19910 0 0 $X=35810 $Y=19660
X73 55 M4_M3_CDNS_7656752519063 $T=44820 19910 0 0 $X=44600 $Y=19660
X74 56 M4_M3_CDNS_7656752519063 $T=50410 19910 0 0 $X=50190 $Y=19660
X75 57 M4_M3_CDNS_7656752519063 $T=53190 19910 0 0 $X=52970 $Y=19660
X76 50 M3_M2_CDNS_7656752519064 $T=9340 19910 0 0 $X=9120 $Y=19660
X77 51 M3_M2_CDNS_7656752519064 $T=18130 19910 0 0 $X=17910 $Y=19660
X78 52 M3_M2_CDNS_7656752519064 $T=23720 19910 0 0 $X=23500 $Y=19660
X79 53 M3_M2_CDNS_7656752519064 $T=26500 19910 0 0 $X=26280 $Y=19660
X80 54 M3_M2_CDNS_7656752519064 $T=36030 19910 0 0 $X=35810 $Y=19660
X81 55 M3_M2_CDNS_7656752519064 $T=44820 19910 0 0 $X=44600 $Y=19660
X82 56 M3_M2_CDNS_7656752519064 $T=50410 19910 0 0 $X=50190 $Y=19660
X83 57 M3_M2_CDNS_7656752519064 $T=53190 19910 0 0 $X=52970 $Y=19660
X84 50 M2_M1_CDNS_7656752519065 $T=9340 19910 0 0 $X=9120 $Y=19660
X85 51 M2_M1_CDNS_7656752519065 $T=18130 19910 0 0 $X=17910 $Y=19660
X86 52 M2_M1_CDNS_7656752519065 $T=23720 19910 0 0 $X=23500 $Y=19660
X87 53 M2_M1_CDNS_7656752519065 $T=26500 19910 0 0 $X=26280 $Y=19660
X88 54 M2_M1_CDNS_7656752519065 $T=36030 19910 0 0 $X=35810 $Y=19660
X89 55 M2_M1_CDNS_7656752519065 $T=44820 19910 0 0 $X=44600 $Y=19660
X90 56 M2_M1_CDNS_7656752519065 $T=50410 19910 0 0 $X=50190 $Y=19660
X91 57 M2_M1_CDNS_7656752519065 $T=53190 19910 0 0 $X=52970 $Y=19660
X92 50 M6_M5_CDNS_7656752519066 $T=9340 19910 0 0 $X=9120 $Y=19660
X93 51 M6_M5_CDNS_7656752519066 $T=18130 19910 0 0 $X=17910 $Y=19660
X94 52 M6_M5_CDNS_7656752519066 $T=23720 19910 0 0 $X=23500 $Y=19660
X95 53 M6_M5_CDNS_7656752519066 $T=26500 19910 0 0 $X=26280 $Y=19660
X96 54 M6_M5_CDNS_7656752519066 $T=36030 19910 0 0 $X=35810 $Y=19660
X97 55 M6_M5_CDNS_7656752519066 $T=44820 19910 0 0 $X=44600 $Y=19660
X98 56 M6_M5_CDNS_7656752519066 $T=50410 19910 0 0 $X=50190 $Y=19660
X99 57 M6_M5_CDNS_7656752519066 $T=53190 19910 0 0 $X=52970 $Y=19660
X100 8 2 6 5 50 66 109 AND $T=3670 21910 0 0 $X=4740 $Y=18810
X101 12 9 6 5 51 70 112 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X102 14 11 6 5 52 73 115 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X103 17 16 6 5 53 80 128 AND $T=32210 21910 1 180 $X=26960 $Y=18810
X104 19 18 6 5 54 82 130 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X105 23 22 6 5 55 86 134 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X106 26 25 6 5 56 89 137 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X107 29 28 6 5 57 94 142 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X108 3 5 6 33 4 106 64 XOR $T=530 18810 1 0 $X=530 $Y=14110
X109 42 5 6 1 33 105 63 XOR $T=640 4700 1 0 $X=640 $Y=0
X110 2 5 6 34 8 108 65 XOR $T=4740 18810 1 0 $X=4740 $Y=14110
X111 43 5 6 7 34 107 67 XOR $T=9740 4700 0 180 $X=6020 $Y=0
X112 44 5 6 10 35 111 69 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X113 9 5 6 35 12 110 68 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X114 45 5 6 13 36 114 72 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X115 11 5 6 36 14 113 71 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X116 46 5 6 15 37 116 74 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X117 16 5 6 37 17 127 79 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X118 18 5 6 38 19 129 81 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X119 47 5 6 20 38 131 83 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X120 48 5 6 21 39 133 85 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X121 22 5 6 39 23 132 84 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X122 49 5 6 24 40 136 88 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X123 25 5 6 40 26 135 87 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X124 58 5 6 27 41 138 90 XOR $T=49650 4700 1 0 $X=49650 $Y=0
X125 28 5 6 41 29 141 93 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X126 30 5 58 31 32 6 92 91 139 163
+ 164 140 HAdder $T=62720 6180 1 90 $X=53760 $Y=6980
X127 37 53 46 5 6 36 52 45 35 51
+ 44 34 43 50 42 59 60 61 62 143
+ 145 144 146 147 148 150 151 152 149 95
+ 96 99 100 98 101 102 97 103 104 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X128 41 57 58 5 6 40 56 49 39 55
+ 48 38 47 54 46 75 76 77 78 153
+ 155 154 156 157 158 160 161 162 159 117
+ 118 121 122 120 123 124 119 125 126 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
M0 109 2 66 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5600 $Y=19150 $dt=0
M1 5 8 109 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5810 $Y=19150 $dt=0
M2 50 66 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=8230 $Y=19140 $dt=0
M3 112 9 70 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=19150 $dt=0
M4 5 12 112 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=19150 $dt=0
M5 51 70 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=19140 $dt=0
M6 115 11 73 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=19150 $dt=0
M7 5 14 115 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=19150 $dt=0
M8 52 73 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=19140 $dt=0
M9 5 80 53 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27560 $Y=19140 $dt=0
M10 128 17 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29980 $Y=19150 $dt=0
M11 80 16 128 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30190 $Y=19150 $dt=0
M12 130 18 82 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=19150 $dt=0
M13 5 19 130 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=19150 $dt=0
M14 54 82 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=19140 $dt=0
M15 134 22 86 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=19150 $dt=0
M16 5 23 134 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=19150 $dt=0
M17 55 86 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=19140 $dt=0
M18 137 25 89 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=19150 $dt=0
M19 5 26 137 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=19150 $dt=0
M20 56 89 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=19140 $dt=0
M21 5 94 57 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=19140 $dt=0
M22 142 29 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=19150 $dt=0
M23 94 28 142 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=19150 $dt=0
M24 6 62 42 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M25 106 3 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=950 $Y=14910 $dt=1
M26 105 42 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=115.144 scb=0.0588049 scc=0.0138331 $X=1060 $Y=800 $dt=1
M27 149 50 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M28 33 4 3 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=1880 $Y=14910 $dt=1
M29 1 33 42 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.854 scb=0.0354545 scc=0.011187 $X=1990 $Y=800 $dt=1
M30 106 64 33 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=2810 $Y=14910 $dt=1
M31 105 63 1 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=2920 $Y=800 $dt=1
M32 6 4 64 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=3740 $Y=14910 $dt=1
M33 6 33 63 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=3850 $Y=800 $dt=1
M34 108 2 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=14910 $dt=1
M35 66 2 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=20590 $dt=1
M36 6 8 66 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=20590 $dt=1
M37 34 8 2 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=14910 $dt=1
M38 67 34 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=6440 $Y=800 $dt=1
M39 108 65 34 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=14910 $dt=1
M40 7 67 107 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=7370 $Y=800 $dt=1
M41 6 8 65 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=14910 $dt=1
M42 50 66 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=8230 $Y=20400 $dt=1
M43 43 34 7 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=8300 $Y=800 $dt=1
M44 6 43 107 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=9230 $Y=800 $dt=1
M45 69 35 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=13880 $Y=800 $dt=1
M46 110 9 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M47 70 9 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=20590 $dt=1
M48 6 12 70 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=20590 $dt=1
M49 10 69 111 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=14810 $Y=800 $dt=1
M50 35 12 9 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M51 44 35 10 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=15740 $Y=800 $dt=1
M52 110 68 35 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M53 6 44 111 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=16670 $Y=800 $dt=1
M54 6 12 68 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M55 51 70 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17020 $Y=20400 $dt=1
M56 72 36 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=19460 $Y=800 $dt=1
M57 113 11 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M58 73 11 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=20590 $dt=1
M59 13 72 114 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=20390 $Y=800 $dt=1
M60 6 14 73 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=20590 $dt=1
M61 36 14 11 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M62 45 36 13 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=21320 $Y=800 $dt=1
M63 113 71 36 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M64 6 45 114 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=22250 $Y=800 $dt=1
M65 6 14 71 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M66 52 73 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22610 $Y=20400 $dt=1
M67 74 37 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=23510 $Y=800 $dt=1
M68 15 74 116 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=24440 $Y=800 $dt=1
M69 46 37 15 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=25370 $Y=800 $dt=1
M70 6 46 116 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=26300 $Y=800 $dt=1
M71 6 78 46 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M72 6 80 53 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27560 $Y=20400 $dt=1
M73 79 17 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M74 159 54 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M75 37 79 127 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M76 16 17 37 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M77 80 17 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29780 $Y=20590 $dt=1
M78 6 16 80 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30190 $Y=20590 $dt=1
M79 6 16 127 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M80 129 18 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M81 82 18 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=20590 $dt=1
M82 6 19 82 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=20590 $dt=1
M83 38 19 18 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M84 83 38 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=33170 $Y=800 $dt=1
M85 129 81 38 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M86 20 83 131 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=34100 $Y=800 $dt=1
M87 6 19 81 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M88 54 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=34920 $Y=20400 $dt=1
M89 47 38 20 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=35030 $Y=800 $dt=1
M90 6 47 131 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35960 $Y=800 $dt=1
M91 85 39 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=40590 $Y=800 $dt=1
M92 132 22 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M93 86 22 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=20590 $dt=1
M94 6 23 86 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=20590 $dt=1
M95 21 85 133 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=41520 $Y=800 $dt=1
M96 39 23 22 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M97 48 39 21 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=42450 $Y=800 $dt=1
M98 132 84 39 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M99 6 48 133 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=43380 $Y=800 $dt=1
M100 6 23 84 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M101 55 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=43710 $Y=20400 $dt=1
M102 88 40 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=46150 $Y=800 $dt=1
M103 135 25 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M104 89 25 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=20590 $dt=1
M105 24 88 136 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=47080 $Y=800 $dt=1
M106 6 26 89 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=20590 $dt=1
M107 40 26 25 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M108 49 40 24 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=48010 $Y=800 $dt=1
M109 135 87 40 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M110 6 49 136 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6675 scb=0.0347689 scc=0.0111862 $X=48940 $Y=800 $dt=1
M111 6 26 87 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M112 56 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=49300 $Y=20400 $dt=1
M113 138 58 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=50070 $Y=800 $dt=1
M114 27 41 58 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51000 $Y=800 $dt=1
M115 138 90 27 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51930 $Y=800 $dt=1
M116 6 41 90 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=52860 $Y=800 $dt=1
M117 6 94 57 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=54210 $Y=20400 $dt=1
M118 93 29 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M119 41 93 141 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M120 164 92 58 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=55830 $Y=11700 $dt=1
M121 6 91 164 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56040 $Y=11700 $dt=1
M122 28 29 41 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M123 94 29 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=20590 $dt=1
M124 6 28 94 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=20590 $dt=1
M125 6 91 163 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56970 $Y=11700 $dt=1
M126 6 28 141 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M127 163 92 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57380 $Y=11700 $dt=1
M128 30 32 163 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57790 $Y=11700 $dt=1
M129 163 31 30 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=58200 $Y=11700 $dt=1
M130 6 31 91 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=59130 $Y=11700 $dt=1
M131 6 32 92 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=60060 $Y=11700 $dt=1
.ends WallaceFinalAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656752519085                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656752519085 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656752519085

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519021                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519021 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656752519021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519022                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519022 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656752519022

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519023                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519023 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656752519023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656752519024                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656752519024 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656752519024

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519025                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519025 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.6986 scb=0.0347897 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656752519025

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519026                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519026 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656752519026

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656752519027                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656752519027 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656752519027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAdder 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=10
X0 8 M2_M1_CDNS_7656752519020 $T=2700 5110 0 90 $X=2570 $Y=5030
X1 9 M2_M1_CDNS_7656752519020 $T=3060 2950 0 90 $X=2930 $Y=2870
X2 9 M2_M1_CDNS_7656752519020 $T=3060 5520 0 90 $X=2930 $Y=5440
X3 5 M2_M1_CDNS_7656752519020 $T=3450 7370 0 90 $X=3320 $Y=7290
X4 3 M2_M1_CDNS_7656752519020 $T=3450 8190 0 90 $X=3320 $Y=8110
X5 5 M2_M1_CDNS_7656752519020 $T=3460 3880 0 90 $X=3330 $Y=3800
X6 3 M2_M1_CDNS_7656752519020 $T=4250 4700 0 90 $X=4120 $Y=4620
X7 10 M2_M1_CDNS_7656752519020 $T=4700 5110 0 90 $X=4570 $Y=5030
X8 10 M2_M1_CDNS_7656752519020 $T=4740 5820 0 90 $X=4610 $Y=5740
X9 8 M2_M1_CDNS_7656752519020 $T=5140 5990 0 90 $X=5010 $Y=5910
X10 8 M2_M1_CDNS_7656752519025 $T=5020 6720 0 90 $X=4890 $Y=6590
X11 10 M1_PO_CDNS_7656752519067 $T=1550 6040 0 90 $X=1430 $Y=5940
X12 5 M1_PO_CDNS_7656752519067 $T=3090 2650 0 90 $X=2970 $Y=2550
X13 5 M1_PO_CDNS_7656752519067 $T=3090 3820 0 90 $X=2970 $Y=3720
X14 5 M1_PO_CDNS_7656752519067 $T=3090 4360 0 90 $X=2970 $Y=4260
X15 6 M1_PO_CDNS_7656752519067 $T=3145 6870 0 90 $X=3025 $Y=6770
X16 9 M1_PO_CDNS_7656752519067 $T=3720 5020 0 90 $X=3600 $Y=4920
X17 8 M1_PO_CDNS_7656752519068 $T=2700 7470 0 90 $X=2450 $Y=7370
X18 6 M1_PO_CDNS_7656752519068 $T=3820 6180 0 90 $X=3570 $Y=6080
X19 3 M1_PO_CDNS_7656752519068 $T=4200 5220 0 90 $X=3950 $Y=5120
X20 3 M1_PO_CDNS_7656752519068 $T=4250 4170 0 90 $X=4000 $Y=4070
X21 10 M1_PO_CDNS_7656752519068 $T=4650 8090 0 90 $X=4400 $Y=7990
X22 8 M1_PO_CDNS_7656752519068 $T=5020 6720 0 90 $X=4770 $Y=6620
X23 8 M2_M1_CDNS_7656752519069 $T=2700 7470 0 90 $X=2450 $Y=7390
X24 6 M2_M1_CDNS_7656752519069 $T=3820 6180 0 90 $X=3570 $Y=6100
X25 3 M2_M1_CDNS_7656752519069 $T=4200 5220 0 90 $X=3950 $Y=5140
X26 3 M2_M1_CDNS_7656752519069 $T=4250 4170 0 90 $X=4000 $Y=4090
X27 10 M2_M1_CDNS_7656752519069 $T=4650 8090 0 90 $X=4400 $Y=8010
X28 9 3 8 1 nmos1v_CDNS_7656752519014 $T=2220 5270 0 90 $X=1780 $Y=5030
X29 10 6 2 1 nmos1v_CDNS_7656752519014 $T=2220 6290 1 270 $X=1780 $Y=5780
X30 3 10 4 1 nmos1v_CDNS_7656752519014 $T=2220 7950 0 90 $X=1780 $Y=7710
X31 5 3 8 1 7 pmos1v_CDNS_7656752519018 $T=5670 4040 0 90 $X=5230 $Y=3620
X32 9 3 10 1 7 pmos1v_CDNS_7656752519018 $T=5670 5360 1 270 $X=5230 $Y=5030
X33 5 8 4 1 7 pmos1v_CDNS_7656752519018 $T=5670 7540 0 90 $X=5230 $Y=7120
X34 7 7 5 9 1 pmos1v_CDNS_7656752519019 $T=5670 3200 1 270 $X=5230 $Y=2690
X35 1 1 5 9 nmos1v_CDNS_7656752519020 $T=2220 3200 1 270 $X=1420 $Y=2690
X36 6 M2_M1_CDNS_7656752519085 $T=3820 2110 0 90 $X=3740 $Y=1860
X37 3 M2_M1_CDNS_7656752519085 $T=4260 2110 0 90 $X=4180 $Y=1860
X38 5 3 10 1 nmos1v_CDNS_7656752519021 $T=2220 4450 0 90 $X=1780 $Y=4210
X39 10 5 3 1 nmos1v_CDNS_7656752519022 $T=2220 4130 1 270 $X=1780 $Y=3620
X40 2 6 10 1 nmos1v_CDNS_7656752519022 $T=2220 6610 0 90 $X=1780 $Y=6250
X41 4 6 8 1 nmos1v_CDNS_7656752519022 $T=2220 7630 1 270 $X=1780 $Y=7120
X42 6 8 2 1 7 pmos1v_CDNS_7656752519023 $T=5670 6700 1 270 $X=5230 $Y=6250
X43 6 10 4 1 7 pmos1v_CDNS_7656752519023 $T=5670 8040 1 270 $X=5230 $Y=7590
X44 8 3 9 1 nmos1v_CDNS_7656752519024 $T=2220 4950 1 270 $X=1780 $Y=4500
X45 8 5 3 1 7 pmos1v_CDNS_7656752519025 $T=5670 4540 1 270 $X=5230 $Y=4090
X46 3 10 9 1 7 pmos1v_CDNS_7656752519026 $T=5670 4860 0 90 $X=5230 $Y=4500
X47 8 6 2 1 7 pmos1v_CDNS_7656752519027 $T=5670 6200 0 90 $X=5230 $Y=5780
M0 4 8 6 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=7540 $dt=0
M1 7 5 9 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5430 $Y=3110 $dt=1
M2 8 3 5 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5430 $Y=4040 $dt=1
M3 9 3 10 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5430 $Y=5270 $dt=1
M4 6 8 2 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=95.6709 scb=0.0347795 scc=0.0111862 $X=5430 $Y=6610 $dt=1
M5 4 8 5 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=99.6807 scb=0.0402027 scc=0.0112574 $X=5430 $Y=7540 $dt=1
.ends FAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y1 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=0
X0 1 M2_M1_CDNS_7656752519028 $T=80 250 0 0 $X=0 $Y=0
X1 2 M2_M1_CDNS_7656752519028 $T=480 250 0 0 $X=400 $Y=0
X2 3 M2_M1_CDNS_7656752519028 $T=880 250 0 0 $X=800 $Y=0
X3 4 M2_M1_CDNS_7656752519028 $T=1280 250 0 0 $X=1200 $Y=0
X4 5 M2_M1_CDNS_7656752519028 $T=1680 250 0 0 $X=1600 $Y=0
X5 6 M2_M1_CDNS_7656752519028 $T=2080 250 0 0 $X=2000 $Y=0
X6 7 M2_M1_CDNS_7656752519028 $T=2480 250 0 0 $X=2400 $Y=0
X7 8 M2_M1_CDNS_7656752519028 $T=2880 250 0 0 $X=2800 $Y=0
.ends MASCO__Y1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y2 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=0
X0 1 M3_M2_CDNS_7656752519027 $T=80 250 0 0 $X=0 $Y=0
X1 2 M3_M2_CDNS_7656752519027 $T=480 250 0 0 $X=400 $Y=0
X2 3 M3_M2_CDNS_7656752519027 $T=880 250 0 0 $X=800 $Y=0
X3 4 M3_M2_CDNS_7656752519027 $T=1280 250 0 0 $X=1200 $Y=0
X4 5 M3_M2_CDNS_7656752519027 $T=1680 250 0 0 $X=1600 $Y=0
X5 6 M3_M2_CDNS_7656752519027 $T=2080 250 0 0 $X=2000 $Y=0
X6 7 M3_M2_CDNS_7656752519027 $T=2480 250 0 0 $X=2400 $Y=0
X7 8 M3_M2_CDNS_7656752519027 $T=2880 250 0 0 $X=2800 $Y=0
.ends MASCO__Y2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceMultiplier                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceMultiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82
** N=210 EP=82 FDC=384
X0 2 M2_M1_CDNS_7656752519020 $T=2220 31930 0 0 $X=2140 $Y=31800
X1 3 M2_M1_CDNS_7656752519020 $T=2220 35820 0 0 $X=2140 $Y=35690
X2 4 M2_M1_CDNS_7656752519020 $T=2220 36470 0 0 $X=2140 $Y=36340
X3 5 M2_M1_CDNS_7656752519020 $T=2220 40360 0 0 $X=2140 $Y=40230
X4 6 M2_M1_CDNS_7656752519020 $T=2220 41010 0 0 $X=2140 $Y=40880
X5 7 M2_M1_CDNS_7656752519020 $T=2220 44900 0 0 $X=2140 $Y=44770
X6 8 M2_M1_CDNS_7656752519020 $T=2220 45540 0 0 $X=2140 $Y=45410
X7 9 M2_M1_CDNS_7656752519020 $T=2220 49430 0 0 $X=2140 $Y=49300
X8 2 M2_M1_CDNS_7656752519020 $T=3380 32500 0 0 $X=3300 $Y=32370
X9 3 M2_M1_CDNS_7656752519020 $T=3380 35240 0 0 $X=3300 $Y=35110
X10 4 M2_M1_CDNS_7656752519020 $T=3380 37040 0 0 $X=3300 $Y=36910
X11 5 M2_M1_CDNS_7656752519020 $T=3380 39780 0 0 $X=3300 $Y=39650
X12 6 M2_M1_CDNS_7656752519020 $T=3380 41580 0 0 $X=3300 $Y=41450
X13 7 M2_M1_CDNS_7656752519020 $T=3380 44320 0 0 $X=3300 $Y=44190
X14 8 M2_M1_CDNS_7656752519020 $T=3380 46120 0 0 $X=3300 $Y=45990
X15 9 M2_M1_CDNS_7656752519020 $T=3380 48860 0 0 $X=3300 $Y=48730
X16 2 M2_M1_CDNS_7656752519020 $T=8590 32500 0 0 $X=8510 $Y=32370
X17 3 M2_M1_CDNS_7656752519020 $T=8590 35240 0 0 $X=8510 $Y=35110
X18 4 M2_M1_CDNS_7656752519020 $T=8590 37040 0 0 $X=8510 $Y=36910
X19 5 M2_M1_CDNS_7656752519020 $T=8590 39780 0 0 $X=8510 $Y=39650
X20 6 M2_M1_CDNS_7656752519020 $T=8590 41580 0 0 $X=8510 $Y=41450
X21 7 M2_M1_CDNS_7656752519020 $T=8590 44320 0 0 $X=8510 $Y=44190
X22 8 M2_M1_CDNS_7656752519020 $T=8590 46120 0 0 $X=8510 $Y=45990
X23 9 M2_M1_CDNS_7656752519020 $T=8590 48860 0 0 $X=8510 $Y=48730
X24 2 M2_M1_CDNS_7656752519020 $T=13610 32500 0 0 $X=13530 $Y=32370
X25 3 M2_M1_CDNS_7656752519020 $T=13610 35240 0 0 $X=13530 $Y=35110
X26 4 M2_M1_CDNS_7656752519020 $T=13610 37040 0 0 $X=13530 $Y=36910
X27 5 M2_M1_CDNS_7656752519020 $T=13610 39780 0 0 $X=13530 $Y=39650
X28 6 M2_M1_CDNS_7656752519020 $T=13610 41580 0 0 $X=13530 $Y=41450
X29 7 M2_M1_CDNS_7656752519020 $T=13610 44320 0 0 $X=13530 $Y=44190
X30 8 M2_M1_CDNS_7656752519020 $T=13610 46120 0 0 $X=13530 $Y=45990
X31 9 M2_M1_CDNS_7656752519020 $T=13610 48860 0 0 $X=13530 $Y=48730
X32 2 M2_M1_CDNS_7656752519020 $T=18740 32500 0 0 $X=18660 $Y=32370
X33 3 M2_M1_CDNS_7656752519020 $T=18740 35240 0 0 $X=18660 $Y=35110
X34 4 M2_M1_CDNS_7656752519020 $T=18740 37040 0 0 $X=18660 $Y=36910
X35 5 M2_M1_CDNS_7656752519020 $T=18740 39780 0 0 $X=18660 $Y=39650
X36 6 M2_M1_CDNS_7656752519020 $T=18740 41580 0 0 $X=18660 $Y=41450
X37 7 M2_M1_CDNS_7656752519020 $T=18740 44320 0 0 $X=18660 $Y=44190
X38 8 M2_M1_CDNS_7656752519020 $T=18740 46120 0 0 $X=18660 $Y=45990
X39 9 M2_M1_CDNS_7656752519020 $T=18740 48860 0 0 $X=18660 $Y=48730
X40 2 M2_M1_CDNS_7656752519020 $T=23810 32500 0 0 $X=23730 $Y=32370
X41 3 M2_M1_CDNS_7656752519020 $T=23810 35240 0 0 $X=23730 $Y=35110
X42 4 M2_M1_CDNS_7656752519020 $T=23810 37040 0 0 $X=23730 $Y=36910
X43 5 M2_M1_CDNS_7656752519020 $T=23810 39780 0 0 $X=23730 $Y=39650
X44 6 M2_M1_CDNS_7656752519020 $T=23810 41580 0 0 $X=23730 $Y=41450
X45 7 M2_M1_CDNS_7656752519020 $T=23810 44320 0 0 $X=23730 $Y=44190
X46 8 M2_M1_CDNS_7656752519020 $T=23810 46120 0 0 $X=23730 $Y=45990
X47 9 M2_M1_CDNS_7656752519020 $T=23810 48860 0 0 $X=23730 $Y=48730
X48 2 M2_M1_CDNS_7656752519020 $T=28690 32500 0 0 $X=28610 $Y=32370
X49 3 M2_M1_CDNS_7656752519020 $T=28690 35240 0 0 $X=28610 $Y=35110
X50 4 M2_M1_CDNS_7656752519020 $T=28690 37040 0 0 $X=28610 $Y=36910
X51 5 M2_M1_CDNS_7656752519020 $T=28690 39780 0 0 $X=28610 $Y=39650
X52 6 M2_M1_CDNS_7656752519020 $T=28690 41580 0 0 $X=28610 $Y=41450
X53 7 M2_M1_CDNS_7656752519020 $T=28690 44320 0 0 $X=28610 $Y=44190
X54 8 M2_M1_CDNS_7656752519020 $T=28690 46120 0 0 $X=28610 $Y=45990
X55 9 M2_M1_CDNS_7656752519020 $T=28690 48860 0 0 $X=28610 $Y=48730
X56 2 M2_M1_CDNS_7656752519020 $T=33890 32500 0 0 $X=33810 $Y=32370
X57 3 M2_M1_CDNS_7656752519020 $T=33890 35240 0 0 $X=33810 $Y=35110
X58 4 M2_M1_CDNS_7656752519020 $T=33890 37040 0 0 $X=33810 $Y=36910
X59 5 M2_M1_CDNS_7656752519020 $T=33890 39780 0 0 $X=33810 $Y=39650
X60 6 M2_M1_CDNS_7656752519020 $T=33890 41580 0 0 $X=33810 $Y=41450
X61 7 M2_M1_CDNS_7656752519020 $T=33890 44320 0 0 $X=33810 $Y=44190
X62 8 M2_M1_CDNS_7656752519020 $T=33890 46120 0 0 $X=33810 $Y=45990
X63 9 M2_M1_CDNS_7656752519020 $T=33890 48860 0 0 $X=33810 $Y=48730
X64 2 M2_M1_CDNS_7656752519020 $T=38920 32500 0 0 $X=38840 $Y=32370
X65 3 M2_M1_CDNS_7656752519020 $T=38920 35240 0 0 $X=38840 $Y=35110
X66 4 M2_M1_CDNS_7656752519020 $T=38920 37040 0 0 $X=38840 $Y=36910
X67 5 M2_M1_CDNS_7656752519020 $T=38920 39780 0 0 $X=38840 $Y=39650
X68 6 M2_M1_CDNS_7656752519020 $T=38920 41580 0 0 $X=38840 $Y=41450
X69 7 M2_M1_CDNS_7656752519020 $T=38920 44320 0 0 $X=38840 $Y=44190
X70 8 M2_M1_CDNS_7656752519020 $T=38920 46120 0 0 $X=38840 $Y=45990
X71 9 M2_M1_CDNS_7656752519020 $T=38920 48860 0 0 $X=38840 $Y=48730
X72 1 M3_M2_CDNS_7656752519027 $T=3380 31230 0 0 $X=3300 $Y=30980
X73 1 M3_M2_CDNS_7656752519027 $T=3380 33140 0 0 $X=3300 $Y=32890
X74 1 M3_M2_CDNS_7656752519027 $T=3380 34600 0 0 $X=3300 $Y=34350
X75 1 M3_M2_CDNS_7656752519027 $T=3380 37680 0 0 $X=3300 $Y=37430
X76 1 M3_M2_CDNS_7656752519027 $T=3380 39140 0 0 $X=3300 $Y=38890
X77 1 M3_M2_CDNS_7656752519027 $T=3380 42220 0 0 $X=3300 $Y=41970
X78 1 M3_M2_CDNS_7656752519027 $T=3380 43680 0 0 $X=3300 $Y=43430
X79 1 M3_M2_CDNS_7656752519027 $T=3380 46750 0 0 $X=3300 $Y=46500
X80 1 M3_M2_CDNS_7656752519027 $T=3380 48210 0 0 $X=3300 $Y=47960
X81 20 M3_M2_CDNS_7656752519027 $T=8570 31230 0 0 $X=8490 $Y=30980
X82 20 M3_M2_CDNS_7656752519027 $T=8570 33140 0 0 $X=8490 $Y=32890
X83 20 M3_M2_CDNS_7656752519027 $T=8570 34600 0 0 $X=8490 $Y=34350
X84 20 M3_M2_CDNS_7656752519027 $T=8570 37680 0 0 $X=8490 $Y=37430
X85 20 M3_M2_CDNS_7656752519027 $T=8570 39140 0 0 $X=8490 $Y=38890
X86 20 M3_M2_CDNS_7656752519027 $T=8570 42220 0 0 $X=8490 $Y=41970
X87 20 M3_M2_CDNS_7656752519027 $T=8570 43680 0 0 $X=8490 $Y=43430
X88 20 M3_M2_CDNS_7656752519027 $T=8570 46750 0 0 $X=8490 $Y=46500
X89 20 M3_M2_CDNS_7656752519027 $T=8570 48210 0 0 $X=8490 $Y=47960
X90 29 M3_M2_CDNS_7656752519027 $T=13600 31060 0 0 $X=13520 $Y=30810
X91 29 M3_M2_CDNS_7656752519027 $T=13600 33140 0 0 $X=13520 $Y=32890
X92 29 M3_M2_CDNS_7656752519027 $T=13600 34600 0 0 $X=13520 $Y=34350
X93 29 M3_M2_CDNS_7656752519027 $T=13600 37680 0 0 $X=13520 $Y=37430
X94 29 M3_M2_CDNS_7656752519027 $T=13600 39140 0 0 $X=13520 $Y=38890
X95 29 M3_M2_CDNS_7656752519027 $T=13600 42220 0 0 $X=13520 $Y=41970
X96 29 M3_M2_CDNS_7656752519027 $T=13600 43680 0 0 $X=13520 $Y=43430
X97 29 M3_M2_CDNS_7656752519027 $T=13600 46750 0 0 $X=13520 $Y=46500
X98 29 M3_M2_CDNS_7656752519027 $T=13600 48210 0 0 $X=13520 $Y=47960
X99 37 M3_M2_CDNS_7656752519027 $T=18750 31230 0 0 $X=18670 $Y=30980
X100 37 M3_M2_CDNS_7656752519027 $T=18750 33140 0 0 $X=18670 $Y=32890
X101 37 M3_M2_CDNS_7656752519027 $T=18750 34600 0 0 $X=18670 $Y=34350
X102 37 M3_M2_CDNS_7656752519027 $T=18750 37680 0 0 $X=18670 $Y=37430
X103 37 M3_M2_CDNS_7656752519027 $T=18750 39140 0 0 $X=18670 $Y=38890
X104 37 M3_M2_CDNS_7656752519027 $T=18750 42220 0 0 $X=18670 $Y=41970
X105 37 M3_M2_CDNS_7656752519027 $T=18750 43680 0 0 $X=18670 $Y=43430
X106 37 M3_M2_CDNS_7656752519027 $T=18750 46750 0 0 $X=18670 $Y=46500
X107 37 M3_M2_CDNS_7656752519027 $T=18750 48210 0 0 $X=18670 $Y=47960
X108 44 M3_M2_CDNS_7656752519027 $T=23840 31230 0 0 $X=23760 $Y=30980
X109 44 M3_M2_CDNS_7656752519027 $T=23840 33140 0 0 $X=23760 $Y=32890
X110 44 M3_M2_CDNS_7656752519027 $T=23840 34600 0 0 $X=23760 $Y=34350
X111 44 M3_M2_CDNS_7656752519027 $T=23840 37680 0 0 $X=23760 $Y=37430
X112 44 M3_M2_CDNS_7656752519027 $T=23840 39140 0 0 $X=23760 $Y=38890
X113 44 M3_M2_CDNS_7656752519027 $T=23840 42220 0 0 $X=23760 $Y=41970
X114 44 M3_M2_CDNS_7656752519027 $T=23840 43680 0 0 $X=23760 $Y=43430
X115 44 M3_M2_CDNS_7656752519027 $T=23840 46750 0 0 $X=23760 $Y=46500
X116 44 M3_M2_CDNS_7656752519027 $T=23840 48210 0 0 $X=23760 $Y=47960
X117 56 M3_M2_CDNS_7656752519027 $T=28730 31230 0 0 $X=28650 $Y=30980
X118 56 M3_M2_CDNS_7656752519027 $T=28730 33140 0 0 $X=28650 $Y=32890
X119 56 M3_M2_CDNS_7656752519027 $T=28730 34600 0 0 $X=28650 $Y=34350
X120 56 M3_M2_CDNS_7656752519027 $T=28730 37680 0 0 $X=28650 $Y=37430
X121 56 M3_M2_CDNS_7656752519027 $T=28730 39140 0 0 $X=28650 $Y=38890
X122 56 M3_M2_CDNS_7656752519027 $T=28730 42220 0 0 $X=28650 $Y=41970
X123 56 M3_M2_CDNS_7656752519027 $T=28730 43680 0 0 $X=28650 $Y=43430
X124 56 M3_M2_CDNS_7656752519027 $T=28730 46750 0 0 $X=28650 $Y=46500
X125 56 M3_M2_CDNS_7656752519027 $T=28730 48210 0 0 $X=28650 $Y=47960
X126 65 M3_M2_CDNS_7656752519027 $T=33970 31230 0 0 $X=33890 $Y=30980
X127 65 M3_M2_CDNS_7656752519027 $T=33970 33140 0 0 $X=33890 $Y=32890
X128 65 M3_M2_CDNS_7656752519027 $T=33970 34600 0 0 $X=33890 $Y=34350
X129 65 M3_M2_CDNS_7656752519027 $T=33970 37680 0 0 $X=33890 $Y=37430
X130 65 M3_M2_CDNS_7656752519027 $T=33970 39140 0 0 $X=33890 $Y=38890
X131 65 M3_M2_CDNS_7656752519027 $T=33970 42220 0 0 $X=33890 $Y=41970
X132 65 M3_M2_CDNS_7656752519027 $T=33970 43680 0 0 $X=33890 $Y=43430
X133 65 M3_M2_CDNS_7656752519027 $T=33970 46750 0 0 $X=33890 $Y=46500
X134 65 M3_M2_CDNS_7656752519027 $T=33970 48210 0 0 $X=33890 $Y=47960
X135 73 M3_M2_CDNS_7656752519027 $T=39020 31230 0 0 $X=38940 $Y=30980
X136 73 M3_M2_CDNS_7656752519027 $T=39020 33140 0 0 $X=38940 $Y=32890
X137 73 M3_M2_CDNS_7656752519027 $T=39020 34600 0 0 $X=38940 $Y=34350
X138 73 M3_M2_CDNS_7656752519027 $T=39020 37680 0 0 $X=38940 $Y=37430
X139 73 M3_M2_CDNS_7656752519027 $T=39020 39140 0 0 $X=38940 $Y=38890
X140 73 M3_M2_CDNS_7656752519027 $T=39020 42220 0 0 $X=38940 $Y=41970
X141 73 M3_M2_CDNS_7656752519027 $T=39020 43680 0 0 $X=38940 $Y=43430
X142 73 M3_M2_CDNS_7656752519027 $T=39020 46750 0 0 $X=38940 $Y=46500
X143 73 M3_M2_CDNS_7656752519027 $T=39020 48210 0 0 $X=38940 $Y=47960
X144 1 M2_M1_CDNS_7656752519028 $T=3380 31230 0 0 $X=3300 $Y=30980
X145 1 M2_M1_CDNS_7656752519028 $T=3380 33140 0 0 $X=3300 $Y=32890
X146 1 M2_M1_CDNS_7656752519028 $T=3380 34600 0 0 $X=3300 $Y=34350
X147 1 M2_M1_CDNS_7656752519028 $T=3380 37680 0 0 $X=3300 $Y=37430
X148 1 M2_M1_CDNS_7656752519028 $T=3380 39140 0 0 $X=3300 $Y=38890
X149 1 M2_M1_CDNS_7656752519028 $T=3380 42220 0 0 $X=3300 $Y=41970
X150 1 M2_M1_CDNS_7656752519028 $T=3380 43680 0 0 $X=3300 $Y=43430
X151 1 M2_M1_CDNS_7656752519028 $T=3380 46750 0 0 $X=3300 $Y=46500
X152 1 M2_M1_CDNS_7656752519028 $T=3380 48210 0 0 $X=3300 $Y=47960
X153 20 M2_M1_CDNS_7656752519028 $T=8570 31230 0 0 $X=8490 $Y=30980
X154 20 M2_M1_CDNS_7656752519028 $T=8570 33140 0 0 $X=8490 $Y=32890
X155 20 M2_M1_CDNS_7656752519028 $T=8570 34600 0 0 $X=8490 $Y=34350
X156 20 M2_M1_CDNS_7656752519028 $T=8570 37680 0 0 $X=8490 $Y=37430
X157 20 M2_M1_CDNS_7656752519028 $T=8570 39140 0 0 $X=8490 $Y=38890
X158 20 M2_M1_CDNS_7656752519028 $T=8570 42220 0 0 $X=8490 $Y=41970
X159 20 M2_M1_CDNS_7656752519028 $T=8570 43680 0 0 $X=8490 $Y=43430
X160 20 M2_M1_CDNS_7656752519028 $T=8570 46750 0 0 $X=8490 $Y=46500
X161 20 M2_M1_CDNS_7656752519028 $T=8570 48210 0 0 $X=8490 $Y=47960
X162 29 M2_M1_CDNS_7656752519028 $T=13600 31060 0 0 $X=13520 $Y=30810
X163 29 M2_M1_CDNS_7656752519028 $T=13600 33140 0 0 $X=13520 $Y=32890
X164 29 M2_M1_CDNS_7656752519028 $T=13600 34600 0 0 $X=13520 $Y=34350
X165 29 M2_M1_CDNS_7656752519028 $T=13600 37680 0 0 $X=13520 $Y=37430
X166 29 M2_M1_CDNS_7656752519028 $T=13600 39140 0 0 $X=13520 $Y=38890
X167 29 M2_M1_CDNS_7656752519028 $T=13600 42220 0 0 $X=13520 $Y=41970
X168 29 M2_M1_CDNS_7656752519028 $T=13600 43680 0 0 $X=13520 $Y=43430
X169 29 M2_M1_CDNS_7656752519028 $T=13600 46750 0 0 $X=13520 $Y=46500
X170 29 M2_M1_CDNS_7656752519028 $T=13600 48210 0 0 $X=13520 $Y=47960
X171 37 M2_M1_CDNS_7656752519028 $T=18750 31230 0 0 $X=18670 $Y=30980
X172 37 M2_M1_CDNS_7656752519028 $T=18750 33140 0 0 $X=18670 $Y=32890
X173 37 M2_M1_CDNS_7656752519028 $T=18750 34600 0 0 $X=18670 $Y=34350
X174 37 M2_M1_CDNS_7656752519028 $T=18750 37680 0 0 $X=18670 $Y=37430
X175 37 M2_M1_CDNS_7656752519028 $T=18750 39140 0 0 $X=18670 $Y=38890
X176 37 M2_M1_CDNS_7656752519028 $T=18750 42220 0 0 $X=18670 $Y=41970
X177 37 M2_M1_CDNS_7656752519028 $T=18750 43680 0 0 $X=18670 $Y=43430
X178 37 M2_M1_CDNS_7656752519028 $T=18750 46750 0 0 $X=18670 $Y=46500
X179 37 M2_M1_CDNS_7656752519028 $T=18750 48210 0 0 $X=18670 $Y=47960
X180 44 M2_M1_CDNS_7656752519028 $T=23840 31230 0 0 $X=23760 $Y=30980
X181 44 M2_M1_CDNS_7656752519028 $T=23840 33140 0 0 $X=23760 $Y=32890
X182 44 M2_M1_CDNS_7656752519028 $T=23840 34600 0 0 $X=23760 $Y=34350
X183 44 M2_M1_CDNS_7656752519028 $T=23840 37680 0 0 $X=23760 $Y=37430
X184 44 M2_M1_CDNS_7656752519028 $T=23840 39140 0 0 $X=23760 $Y=38890
X185 44 M2_M1_CDNS_7656752519028 $T=23840 42220 0 0 $X=23760 $Y=41970
X186 44 M2_M1_CDNS_7656752519028 $T=23840 43680 0 0 $X=23760 $Y=43430
X187 44 M2_M1_CDNS_7656752519028 $T=23840 46750 0 0 $X=23760 $Y=46500
X188 44 M2_M1_CDNS_7656752519028 $T=23840 48210 0 0 $X=23760 $Y=47960
X189 56 M2_M1_CDNS_7656752519028 $T=28730 31230 0 0 $X=28650 $Y=30980
X190 56 M2_M1_CDNS_7656752519028 $T=28730 33140 0 0 $X=28650 $Y=32890
X191 56 M2_M1_CDNS_7656752519028 $T=28730 34600 0 0 $X=28650 $Y=34350
X192 56 M2_M1_CDNS_7656752519028 $T=28730 37680 0 0 $X=28650 $Y=37430
X193 56 M2_M1_CDNS_7656752519028 $T=28730 39140 0 0 $X=28650 $Y=38890
X194 56 M2_M1_CDNS_7656752519028 $T=28730 42220 0 0 $X=28650 $Y=41970
X195 56 M2_M1_CDNS_7656752519028 $T=28730 43680 0 0 $X=28650 $Y=43430
X196 56 M2_M1_CDNS_7656752519028 $T=28730 46750 0 0 $X=28650 $Y=46500
X197 56 M2_M1_CDNS_7656752519028 $T=28730 48210 0 0 $X=28650 $Y=47960
X198 65 M2_M1_CDNS_7656752519028 $T=33970 31230 0 0 $X=33890 $Y=30980
X199 65 M2_M1_CDNS_7656752519028 $T=33970 33140 0 0 $X=33890 $Y=32890
X200 65 M2_M1_CDNS_7656752519028 $T=33970 34600 0 0 $X=33890 $Y=34350
X201 65 M2_M1_CDNS_7656752519028 $T=33970 37680 0 0 $X=33890 $Y=37430
X202 65 M2_M1_CDNS_7656752519028 $T=33970 39140 0 0 $X=33890 $Y=38890
X203 65 M2_M1_CDNS_7656752519028 $T=33970 42220 0 0 $X=33890 $Y=41970
X204 65 M2_M1_CDNS_7656752519028 $T=33970 43680 0 0 $X=33890 $Y=43430
X205 65 M2_M1_CDNS_7656752519028 $T=33970 46750 0 0 $X=33890 $Y=46500
X206 65 M2_M1_CDNS_7656752519028 $T=33970 48210 0 0 $X=33890 $Y=47960
X207 73 M2_M1_CDNS_7656752519028 $T=39020 31230 0 0 $X=38940 $Y=30980
X208 73 M2_M1_CDNS_7656752519028 $T=39020 33140 0 0 $X=38940 $Y=32890
X209 73 M2_M1_CDNS_7656752519028 $T=39020 34600 0 0 $X=38940 $Y=34350
X210 73 M2_M1_CDNS_7656752519028 $T=39020 37680 0 0 $X=38940 $Y=37430
X211 73 M2_M1_CDNS_7656752519028 $T=39020 39140 0 0 $X=38940 $Y=38890
X212 73 M2_M1_CDNS_7656752519028 $T=39020 42220 0 0 $X=38940 $Y=41970
X213 73 M2_M1_CDNS_7656752519028 $T=39020 43680 0 0 $X=38940 $Y=43430
X214 73 M2_M1_CDNS_7656752519028 $T=39020 46750 0 0 $X=38940 $Y=46500
X215 73 M2_M1_CDNS_7656752519028 $T=39020 48210 0 0 $X=38940 $Y=47960
X216 1 2 10 16 17 90 154 AND $T=2730 30830 1 0 $X=3800 $Y=31540
X217 1 3 10 16 18 89 153 AND $T=2730 36910 0 0 $X=3800 $Y=33810
X218 1 4 10 16 19 88 152 AND $T=2730 35370 1 0 $X=3800 $Y=36080
X219 1 5 10 16 11 87 151 AND $T=2730 41450 0 0 $X=3800 $Y=38350
X220 1 6 10 16 12 86 150 AND $T=2730 39910 1 0 $X=3800 $Y=40620
X221 1 7 10 16 13 85 149 AND $T=2730 45990 0 0 $X=3800 $Y=42890
X222 1 8 10 16 14 84 148 AND $T=2730 44450 1 0 $X=3800 $Y=45160
X223 1 9 10 16 15 83 147 AND $T=2730 50530 0 0 $X=3800 $Y=47430
X224 20 2 10 16 24 98 162 AND $T=7940 30820 1 0 $X=9010 $Y=31530
X225 20 3 10 16 25 97 161 AND $T=7940 36900 0 0 $X=9010 $Y=33800
X226 20 4 10 16 26 96 160 AND $T=7940 35370 1 0 $X=9010 $Y=36080
X227 20 5 10 16 27 95 159 AND $T=7940 41450 0 0 $X=9010 $Y=38350
X228 20 6 10 16 28 94 158 AND $T=7940 39910 1 0 $X=9010 $Y=40620
X229 20 7 10 16 21 93 157 AND $T=7940 45990 0 0 $X=9010 $Y=42890
X230 20 8 10 16 22 92 156 AND $T=7940 44450 1 0 $X=9010 $Y=45160
X231 20 9 10 16 23 91 155 AND $T=7940 50530 0 0 $X=9010 $Y=47430
X232 29 2 10 16 38 106 170 AND $T=12940 30820 1 0 $X=14010 $Y=31530
X233 29 3 10 16 31 105 169 AND $T=12940 36900 0 0 $X=14010 $Y=33800
X234 29 4 10 16 32 104 168 AND $T=12940 35370 1 0 $X=14010 $Y=36080
X235 29 5 10 16 33 103 167 AND $T=12940 41450 0 0 $X=14010 $Y=38350
X236 29 6 10 16 34 102 166 AND $T=12940 39910 1 0 $X=14010 $Y=40620
X237 29 7 10 16 35 101 165 AND $T=12940 45990 0 0 $X=14010 $Y=42890
X238 29 8 10 16 36 100 164 AND $T=12940 44450 1 0 $X=14010 $Y=45160
X239 29 9 10 16 30 99 163 AND $T=12940 50530 0 0 $X=14010 $Y=47430
X240 37 2 10 16 45 114 178 AND $T=18070 30820 1 0 $X=19140 $Y=31530
X241 37 3 10 16 46 113 177 AND $T=18070 36900 0 0 $X=19140 $Y=33800
X242 37 4 10 16 47 112 176 AND $T=18070 35370 1 0 $X=19140 $Y=36080
X243 37 5 10 16 39 111 175 AND $T=18070 41450 0 0 $X=19140 $Y=38350
X244 37 6 10 16 40 110 174 AND $T=18070 39910 1 0 $X=19140 $Y=40620
X245 37 7 10 16 41 109 173 AND $T=18070 45990 0 0 $X=19140 $Y=42890
X246 37 8 10 16 42 108 172 AND $T=18070 44450 1 0 $X=19140 $Y=45160
X247 37 9 10 16 43 107 171 AND $T=18070 50530 0 0 $X=19140 $Y=47430
X248 44 2 10 16 52 122 186 AND $T=23140 30820 1 0 $X=24210 $Y=31530
X249 44 3 10 16 53 121 185 AND $T=23140 36900 0 0 $X=24210 $Y=33800
X250 44 4 10 16 54 120 184 AND $T=23140 35370 1 0 $X=24210 $Y=36080
X251 44 5 10 16 55 119 183 AND $T=23140 41450 0 0 $X=24210 $Y=38350
X252 44 6 10 16 48 118 182 AND $T=23140 39910 1 0 $X=24210 $Y=40620
X253 44 7 10 16 49 117 181 AND $T=23140 45990 0 0 $X=24210 $Y=42890
X254 44 8 10 16 50 116 180 AND $T=23140 44450 1 0 $X=24210 $Y=45160
X255 44 9 10 16 51 115 179 AND $T=23140 50530 0 0 $X=24210 $Y=47430
X256 56 2 10 16 60 130 194 AND $T=28010 30820 1 0 $X=29080 $Y=31530
X257 56 3 10 16 61 129 193 AND $T=28010 36900 0 0 $X=29080 $Y=33800
X258 56 4 10 16 62 128 192 AND $T=28010 35370 1 0 $X=29080 $Y=36080
X259 56 5 10 16 63 127 191 AND $T=28010 41450 0 0 $X=29080 $Y=38350
X260 56 6 10 16 64 126 190 AND $T=28010 39910 1 0 $X=29080 $Y=40620
X261 56 7 10 16 57 125 189 AND $T=28010 45990 0 0 $X=29080 $Y=42890
X262 56 8 10 16 58 124 188 AND $T=28010 44450 1 0 $X=29080 $Y=45160
X263 56 9 10 16 59 123 187 AND $T=28010 50530 0 0 $X=29080 $Y=47430
X264 65 2 10 16 74 138 202 AND $T=33230 30830 1 0 $X=34300 $Y=31540
X265 65 3 10 16 67 137 201 AND $T=33230 36900 0 0 $X=34300 $Y=33800
X266 65 4 10 16 68 136 200 AND $T=33230 35370 1 0 $X=34300 $Y=36080
X267 65 5 10 16 69 135 199 AND $T=33230 41450 0 0 $X=34300 $Y=38350
X268 65 6 10 16 70 134 198 AND $T=33230 39910 1 0 $X=34300 $Y=40620
X269 65 7 10 16 71 133 197 AND $T=33230 45990 0 0 $X=34300 $Y=42890
X270 65 8 10 16 72 132 196 AND $T=33230 44450 1 0 $X=34300 $Y=45160
X271 65 9 10 16 66 131 195 AND $T=33230 50530 0 0 $X=34300 $Y=47430
X272 73 2 10 16 80 146 210 AND $T=38250 30830 1 0 $X=39320 $Y=31540
X273 73 3 10 16 81 145 209 AND $T=38250 36910 0 0 $X=39320 $Y=33810
X274 73 4 10 16 82 144 208 AND $T=38250 35370 1 0 $X=39320 $Y=36080
X275 73 5 10 16 75 143 207 AND $T=38250 41450 0 0 $X=39320 $Y=38350
X276 73 6 10 16 76 142 206 AND $T=38250 39910 1 0 $X=39320 $Y=40620
X277 73 7 10 16 77 141 205 AND $T=38250 45990 0 0 $X=39320 $Y=42890
X278 73 8 10 16 78 140 204 AND $T=38250 44450 1 0 $X=39320 $Y=45160
X279 73 9 10 16 79 139 203 AND $T=38250 50530 0 0 $X=39320 $Y=47430
X280 15 14 13 12 11 19 18 17 MASCO__Y1 $T=4320 31030 0 0 $X=4320 $Y=31030
X281 23 22 21 28 27 26 25 24 MASCO__Y1 $T=9530 31030 0 0 $X=9530 $Y=31030
X282 30 36 35 34 33 32 31 38 MASCO__Y1 $T=14515 31030 0 0 $X=14515 $Y=31030
X283 43 42 41 40 39 47 46 45 MASCO__Y1 $T=19655 31030 0 0 $X=19655 $Y=31030
X284 51 50 49 48 55 54 53 52 MASCO__Y1 $T=24735 31030 0 0 $X=24735 $Y=31030
X285 59 58 57 64 63 62 61 60 MASCO__Y1 $T=29595 31030 0 0 $X=29595 $Y=31030
X286 66 72 71 70 69 68 67 74 MASCO__Y1 $T=34815 31030 0 0 $X=34815 $Y=31030
X287 79 78 77 76 75 82 81 80 MASCO__Y1 $T=39840 31030 0 0 $X=39840 $Y=31030
X288 15 14 13 12 11 19 18 17 MASCO__Y2 $T=4320 31030 0 0 $X=4320 $Y=31030
X289 23 22 21 28 27 26 25 24 MASCO__Y2 $T=9530 31030 0 0 $X=9530 $Y=31030
X290 30 36 35 34 33 32 31 38 MASCO__Y2 $T=14515 31030 0 0 $X=14515 $Y=31030
X291 43 42 41 40 39 47 46 45 MASCO__Y2 $T=19655 31030 0 0 $X=19655 $Y=31030
X292 51 50 49 48 55 54 53 52 MASCO__Y2 $T=24735 31030 0 0 $X=24735 $Y=31030
X293 59 58 57 64 63 62 61 60 MASCO__Y2 $T=29595 31030 0 0 $X=29595 $Y=31030
X294 66 72 71 70 69 68 67 74 MASCO__Y2 $T=34815 31030 0 0 $X=34815 $Y=31030
X295 79 78 77 76 75 82 81 80 MASCO__Y2 $T=39840 31030 0 0 $X=39840 $Y=31030
M0 154 2 90 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=33350 $dt=0
M1 153 3 89 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=34150 $dt=0
M2 152 4 88 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=37890 $dt=0
M3 151 5 87 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=38690 $dt=0
M4 150 6 86 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=42430 $dt=0
M5 149 7 85 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=43230 $dt=0
M6 148 8 84 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=46970 $dt=0
M7 147 9 83 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=47770 $dt=0
M8 16 1 154 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=33350 $dt=0
M9 16 1 153 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=34150 $dt=0
M10 16 1 152 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=37890 $dt=0
M11 16 1 151 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=38690 $dt=0
M12 16 1 150 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=42430 $dt=0
M13 16 1 149 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=43230 $dt=0
M14 16 1 148 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=46970 $dt=0
M15 16 1 147 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=47770 $dt=0
M16 17 90 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=33360 $dt=0
M17 18 89 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=34140 $dt=0
M18 19 88 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=37900 $dt=0
M19 11 87 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=38680 $dt=0
M20 12 86 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=42440 $dt=0
M21 13 85 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=43220 $dt=0
M22 14 84 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=46980 $dt=0
M23 15 83 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=47760 $dt=0
M24 162 2 98 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=33340 $dt=0
M25 161 3 97 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=34140 $dt=0
M26 160 4 96 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=37890 $dt=0
M27 159 5 95 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=38690 $dt=0
M28 158 6 94 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=42430 $dt=0
M29 157 7 93 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=43230 $dt=0
M30 156 8 92 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=46970 $dt=0
M31 155 9 91 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=47770 $dt=0
M32 16 20 162 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=33340 $dt=0
M33 16 20 161 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=34140 $dt=0
M34 16 20 160 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=37890 $dt=0
M35 16 20 159 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=38690 $dt=0
M36 16 20 158 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=42430 $dt=0
M37 16 20 157 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=43230 $dt=0
M38 16 20 156 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=46970 $dt=0
M39 16 20 155 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=47770 $dt=0
M40 24 98 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=33350 $dt=0
M41 25 97 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=34130 $dt=0
M42 26 96 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=37900 $dt=0
M43 27 95 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=38680 $dt=0
M44 28 94 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=42440 $dt=0
M45 21 93 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=43220 $dt=0
M46 22 92 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=46980 $dt=0
M47 23 91 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=47760 $dt=0
M48 170 2 106 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=33340 $dt=0
M49 169 3 105 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=34140 $dt=0
M50 168 4 104 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=37890 $dt=0
M51 167 5 103 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=38690 $dt=0
M52 166 6 102 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=42430 $dt=0
M53 165 7 101 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=43230 $dt=0
M54 164 8 100 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=46970 $dt=0
M55 163 9 99 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=47770 $dt=0
M56 16 29 170 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=33340 $dt=0
M57 16 29 169 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=34140 $dt=0
M58 16 29 168 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=37890 $dt=0
M59 16 29 167 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=38690 $dt=0
M60 16 29 166 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=42430 $dt=0
M61 16 29 165 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=43230 $dt=0
M62 16 29 164 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=46970 $dt=0
M63 16 29 163 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=47770 $dt=0
M64 38 106 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=33350 $dt=0
M65 31 105 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=34130 $dt=0
M66 32 104 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=37900 $dt=0
M67 33 103 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=38680 $dt=0
M68 34 102 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=42440 $dt=0
M69 35 101 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=43220 $dt=0
M70 36 100 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=46980 $dt=0
M71 30 99 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=47760 $dt=0
M72 178 2 114 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=33340 $dt=0
M73 177 3 113 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=34140 $dt=0
M74 176 4 112 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=37890 $dt=0
M75 175 5 111 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=38690 $dt=0
M76 174 6 110 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=42430 $dt=0
M77 173 7 109 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=43230 $dt=0
M78 172 8 108 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=46970 $dt=0
M79 171 9 107 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=47770 $dt=0
M80 16 37 178 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=33340 $dt=0
M81 16 37 177 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=34140 $dt=0
M82 16 37 176 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=37890 $dt=0
M83 16 37 175 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=38690 $dt=0
M84 16 37 174 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=42430 $dt=0
M85 16 37 173 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=43230 $dt=0
M86 16 37 172 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=46970 $dt=0
M87 16 37 171 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=47770 $dt=0
M88 45 114 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=33350 $dt=0
M89 46 113 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=34130 $dt=0
M90 47 112 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=37900 $dt=0
M91 39 111 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=38680 $dt=0
M92 40 110 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=42440 $dt=0
M93 41 109 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=43220 $dt=0
M94 42 108 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=46980 $dt=0
M95 43 107 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=47760 $dt=0
M96 186 2 122 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=33340 $dt=0
M97 185 3 121 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=34140 $dt=0
M98 184 4 120 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=37890 $dt=0
M99 183 5 119 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=38690 $dt=0
M100 182 6 118 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=42430 $dt=0
M101 181 7 117 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=43230 $dt=0
M102 180 8 116 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=46970 $dt=0
M103 179 9 115 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=47770 $dt=0
M104 16 44 186 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=33340 $dt=0
M105 16 44 185 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=34140 $dt=0
M106 16 44 184 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=37890 $dt=0
M107 16 44 183 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=38690 $dt=0
M108 16 44 182 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=42430 $dt=0
M109 16 44 181 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=43230 $dt=0
M110 16 44 180 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=46970 $dt=0
M111 16 44 179 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=47770 $dt=0
M112 52 122 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=33350 $dt=0
M113 53 121 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=34130 $dt=0
M114 54 120 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=37900 $dt=0
M115 55 119 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=38680 $dt=0
M116 48 118 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=42440 $dt=0
M117 49 117 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=43220 $dt=0
M118 50 116 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=46980 $dt=0
M119 51 115 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=47760 $dt=0
M120 194 2 130 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=33340 $dt=0
M121 193 3 129 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=34140 $dt=0
M122 192 4 128 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=37890 $dt=0
M123 191 5 127 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=38690 $dt=0
M124 190 6 126 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=42430 $dt=0
M125 189 7 125 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=43230 $dt=0
M126 188 8 124 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=46970 $dt=0
M127 187 9 123 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=47770 $dt=0
M128 16 56 194 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=33340 $dt=0
M129 16 56 193 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=34140 $dt=0
M130 16 56 192 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=37890 $dt=0
M131 16 56 191 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=38690 $dt=0
M132 16 56 190 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=42430 $dt=0
M133 16 56 189 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=43230 $dt=0
M134 16 56 188 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=46970 $dt=0
M135 16 56 187 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=47770 $dt=0
M136 60 130 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=33350 $dt=0
M137 61 129 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=34130 $dt=0
M138 62 128 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=37900 $dt=0
M139 63 127 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=38680 $dt=0
M140 64 126 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=42440 $dt=0
M141 57 125 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=43220 $dt=0
M142 58 124 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=46980 $dt=0
M143 59 123 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=47760 $dt=0
M144 202 2 138 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=33350 $dt=0
M145 201 3 137 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=34140 $dt=0
M146 200 4 136 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=37890 $dt=0
M147 199 5 135 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=38690 $dt=0
M148 198 6 134 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=42430 $dt=0
M149 197 7 133 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=43230 $dt=0
M150 196 8 132 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=46970 $dt=0
M151 195 9 131 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=47770 $dt=0
M152 16 65 202 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=33350 $dt=0
M153 16 65 201 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=34140 $dt=0
M154 16 65 200 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=37890 $dt=0
M155 16 65 199 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=38690 $dt=0
M156 16 65 198 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=42430 $dt=0
M157 16 65 197 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=43230 $dt=0
M158 16 65 196 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=46970 $dt=0
M159 16 65 195 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=47770 $dt=0
M160 74 138 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=33360 $dt=0
M161 67 137 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=34130 $dt=0
M162 68 136 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=37900 $dt=0
M163 69 135 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=38680 $dt=0
M164 70 134 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=42440 $dt=0
M165 71 133 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=43220 $dt=0
M166 72 132 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=46980 $dt=0
M167 66 131 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=47760 $dt=0
M168 210 2 146 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=33350 $dt=0
M169 209 3 145 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=34150 $dt=0
M170 208 4 144 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=37890 $dt=0
M171 207 5 143 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=38690 $dt=0
M172 206 6 142 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=42430 $dt=0
M173 205 7 141 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=43230 $dt=0
M174 204 8 140 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=46970 $dt=0
M175 203 9 139 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=47770 $dt=0
M176 16 73 210 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=33350 $dt=0
M177 16 73 209 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=34150 $dt=0
M178 16 73 208 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=37890 $dt=0
M179 16 73 207 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=38690 $dt=0
M180 16 73 206 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=42430 $dt=0
M181 16 73 205 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=43230 $dt=0
M182 16 73 204 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=46970 $dt=0
M183 16 73 203 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=47770 $dt=0
M184 80 146 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=33360 $dt=0
M185 81 145 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=34140 $dt=0
M186 82 144 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=37900 $dt=0
M187 75 143 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=38680 $dt=0
M188 76 142 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=42440 $dt=0
M189 77 141 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=43220 $dt=0
M190 78 140 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=46980 $dt=0
M191 79 139 16 16 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=47760 $dt=0
M192 90 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=31910 $dt=1
M193 89 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=35590 $dt=1
M194 88 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=36450 $dt=1
M195 87 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40130 $dt=1
M196 86 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40990 $dt=1
M197 85 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=44670 $dt=1
M198 84 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=45530 $dt=1
M199 83 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=49210 $dt=1
M200 10 1 90 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=31910 $dt=1
M201 10 1 89 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=35590 $dt=1
M202 10 1 88 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=36450 $dt=1
M203 10 1 87 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40130 $dt=1
M204 10 1 86 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40990 $dt=1
M205 10 1 85 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=44670 $dt=1
M206 10 1 84 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=45530 $dt=1
M207 10 1 83 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=49210 $dt=1
M208 17 90 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=31860 $dt=1
M209 18 89 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=35400 $dt=1
M210 19 88 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=36400 $dt=1
M211 11 87 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=39940 $dt=1
M212 12 86 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=40940 $dt=1
M213 13 85 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=44480 $dt=1
M214 14 84 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=45480 $dt=1
M215 15 83 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=49020 $dt=1
M216 98 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=31900 $dt=1
M217 97 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=35580 $dt=1
M218 96 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=36450 $dt=1
M219 95 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40130 $dt=1
M220 94 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40990 $dt=1
M221 93 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=44670 $dt=1
M222 92 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=45530 $dt=1
M223 91 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=49210 $dt=1
M224 10 20 98 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=31900 $dt=1
M225 10 20 97 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=35580 $dt=1
M226 10 20 96 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=36450 $dt=1
M227 10 20 95 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40130 $dt=1
M228 10 20 94 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40990 $dt=1
M229 10 20 93 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=44670 $dt=1
M230 10 20 92 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=45530 $dt=1
M231 10 20 91 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=49210 $dt=1
M232 24 98 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=31850 $dt=1
M233 25 97 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=35390 $dt=1
M234 26 96 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=36400 $dt=1
M235 27 95 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=39940 $dt=1
M236 28 94 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=40940 $dt=1
M237 21 93 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=44480 $dt=1
M238 22 92 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=45480 $dt=1
M239 23 91 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=49020 $dt=1
M240 106 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=31900 $dt=1
M241 105 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=35580 $dt=1
M242 104 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=36450 $dt=1
M243 103 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40130 $dt=1
M244 102 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40990 $dt=1
M245 101 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=44670 $dt=1
M246 100 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=45530 $dt=1
M247 99 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=49210 $dt=1
M248 10 29 106 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=31900 $dt=1
M249 10 29 105 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=35580 $dt=1
M250 10 29 104 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=36450 $dt=1
M251 10 29 103 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40130 $dt=1
M252 10 29 102 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40990 $dt=1
M253 10 29 101 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=44670 $dt=1
M254 10 29 100 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=45530 $dt=1
M255 10 29 99 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=49210 $dt=1
M256 38 106 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=31850 $dt=1
M257 31 105 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=35390 $dt=1
M258 32 104 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=36400 $dt=1
M259 33 103 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=39940 $dt=1
M260 34 102 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=40940 $dt=1
M261 35 101 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=44480 $dt=1
M262 36 100 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=45480 $dt=1
M263 30 99 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=49020 $dt=1
M264 114 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=31900 $dt=1
M265 113 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=35580 $dt=1
M266 112 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=36450 $dt=1
M267 111 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40130 $dt=1
M268 110 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40990 $dt=1
M269 109 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=44670 $dt=1
M270 108 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=45530 $dt=1
M271 107 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=49210 $dt=1
M272 10 37 114 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=31900 $dt=1
M273 10 37 113 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=35580 $dt=1
M274 10 37 112 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=36450 $dt=1
M275 10 37 111 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40130 $dt=1
M276 10 37 110 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40990 $dt=1
M277 10 37 109 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=44670 $dt=1
M278 10 37 108 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=45530 $dt=1
M279 10 37 107 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=49210 $dt=1
M280 45 114 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=31850 $dt=1
M281 46 113 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=35390 $dt=1
M282 47 112 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=36400 $dt=1
M283 39 111 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=39940 $dt=1
M284 40 110 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=40940 $dt=1
M285 41 109 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=44480 $dt=1
M286 42 108 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=45480 $dt=1
M287 43 107 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=49020 $dt=1
M288 122 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=31900 $dt=1
M289 121 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=35580 $dt=1
M290 120 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=36450 $dt=1
M291 119 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40130 $dt=1
M292 118 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40990 $dt=1
M293 117 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=44670 $dt=1
M294 116 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=45530 $dt=1
M295 115 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=49210 $dt=1
M296 10 44 122 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=31900 $dt=1
M297 10 44 121 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=35580 $dt=1
M298 10 44 120 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=36450 $dt=1
M299 10 44 119 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40130 $dt=1
M300 10 44 118 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40990 $dt=1
M301 10 44 117 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=44670 $dt=1
M302 10 44 116 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=45530 $dt=1
M303 10 44 115 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=49210 $dt=1
M304 52 122 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=31850 $dt=1
M305 53 121 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=35390 $dt=1
M306 54 120 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=36400 $dt=1
M307 55 119 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=39940 $dt=1
M308 48 118 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=40940 $dt=1
M309 49 117 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=44480 $dt=1
M310 50 116 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=45480 $dt=1
M311 51 115 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=49020 $dt=1
M312 130 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=31900 $dt=1
M313 129 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=35580 $dt=1
M314 128 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=36450 $dt=1
M315 127 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40130 $dt=1
M316 126 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40990 $dt=1
M317 125 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=44670 $dt=1
M318 124 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=45530 $dt=1
M319 123 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=49210 $dt=1
M320 10 56 130 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=31900 $dt=1
M321 10 56 129 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=35580 $dt=1
M322 10 56 128 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=36450 $dt=1
M323 10 56 127 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40130 $dt=1
M324 10 56 126 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40990 $dt=1
M325 10 56 125 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=44670 $dt=1
M326 10 56 124 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=45530 $dt=1
M327 10 56 123 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=49210 $dt=1
M328 60 130 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=31850 $dt=1
M329 61 129 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=35390 $dt=1
M330 62 128 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=36400 $dt=1
M331 63 127 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=39940 $dt=1
M332 64 126 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=40940 $dt=1
M333 57 125 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=44480 $dt=1
M334 58 124 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=45480 $dt=1
M335 59 123 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=49020 $dt=1
M336 138 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=31910 $dt=1
M337 137 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=35580 $dt=1
M338 136 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=36450 $dt=1
M339 135 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40130 $dt=1
M340 134 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40990 $dt=1
M341 133 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=44670 $dt=1
M342 132 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=45530 $dt=1
M343 131 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=49210 $dt=1
M344 10 65 138 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=31910 $dt=1
M345 10 65 137 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=35580 $dt=1
M346 10 65 136 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=36450 $dt=1
M347 10 65 135 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40130 $dt=1
M348 10 65 134 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40990 $dt=1
M349 10 65 133 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=44670 $dt=1
M350 10 65 132 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=45530 $dt=1
M351 10 65 131 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=49210 $dt=1
M352 74 138 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=31860 $dt=1
M353 67 137 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=35390 $dt=1
M354 68 136 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=36400 $dt=1
M355 69 135 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=39940 $dt=1
M356 70 134 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=40940 $dt=1
M357 71 133 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=44480 $dt=1
M358 72 132 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=45480 $dt=1
M359 66 131 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=49020 $dt=1
M360 146 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=31910 $dt=1
M361 145 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=35590 $dt=1
M362 144 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=36450 $dt=1
M363 143 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40130 $dt=1
M364 142 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40990 $dt=1
M365 141 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=44670 $dt=1
M366 140 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=45530 $dt=1
M367 139 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=49210 $dt=1
M368 10 73 146 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=31910 $dt=1
M369 10 73 145 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=35590 $dt=1
M370 10 73 144 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=36450 $dt=1
M371 10 73 143 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40130 $dt=1
M372 10 73 142 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40990 $dt=1
M373 10 73 141 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=44670 $dt=1
M374 10 73 140 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=45530 $dt=1
M375 10 73 139 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=49210 $dt=1
M376 80 146 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=31860 $dt=1
M377 81 145 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=35400 $dt=1
M378 82 144 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=36400 $dt=1
M379 75 143 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=39940 $dt=1
M380 76 142 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=40940 $dt=1
M381 77 141 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=44480 $dt=1
M382 78 140 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=45480 $dt=1
M383 79 139 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=49020 $dt=1
.ends WallaceMultiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: Diver                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt Diver 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
X0 2 M1_PO_CDNS_7656752519067 $T=1260 -2440 0 0 $X=1160 $Y=-2560
X1 5 M1_PO_CDNS_7656752519067 $T=2200 -2440 0 0 $X=2100 $Y=-2560
X2 3 3 2 5 1 pmos1v_CDNS_765675251906 $T=1340 -2060 0 0 $X=920 $Y=-2260
X3 3 3 5 4 1 pmos1v_CDNS_765675251906 $T=2270 -2060 0 0 $X=1850 $Y=-2260
X4 1 1 2 5 nmos1v_CDNS_765675251907 $T=1340 -3070 0 0 $X=920 $Y=-3630
X5 1 1 5 4 nmos1v_CDNS_765675251907 $T=2270 -3070 0 0 $X=1850 $Y=-3630
.ends Diver

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MAC                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MAC 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99
** N=291 EP=99 FDC=570
X0 52 M4_M3_CDNS_765675251904 $T=57860 9670 0 90 $X=57730 $Y=9590
X1 5 M2_M1_CDNS_765675251909 $T=9840 3330 0 0 $X=9760 $Y=3080
X2 53 M4_M3_CDNS_7656752519010 $T=150 23850 0 0 $X=70 $Y=23600
X3 54 M4_M3_CDNS_7656752519010 $T=5940 23850 0 0 $X=5860 $Y=23600
X4 55 M4_M3_CDNS_7656752519010 $T=16170 2650 0 0 $X=16090 $Y=2400
X5 56 M4_M3_CDNS_7656752519010 $T=16170 23850 0 0 $X=16090 $Y=23600
X6 57 M4_M3_CDNS_7656752519010 $T=21750 2650 0 0 $X=21670 $Y=2400
X7 58 M4_M3_CDNS_7656752519010 $T=21750 23850 0 0 $X=21670 $Y=23600
X8 59 M4_M3_CDNS_7656752519010 $T=26890 2650 0 0 $X=26810 $Y=2400
X9 60 M4_M3_CDNS_7656752519010 $T=26890 23850 0 0 $X=26810 $Y=23600
X10 61 M4_M3_CDNS_7656752519010 $T=32670 2650 0 0 $X=32590 $Y=2400
X11 62 M4_M3_CDNS_7656752519010 $T=32670 23850 0 0 $X=32590 $Y=23600
X12 63 M4_M3_CDNS_7656752519010 $T=40090 2650 0 0 $X=40010 $Y=2400
X13 64 M4_M3_CDNS_7656752519010 $T=40090 23850 0 0 $X=40010 $Y=23600
X14 65 M4_M3_CDNS_7656752519010 $T=48440 2650 0 0 $X=48360 $Y=2400
X15 66 M4_M3_CDNS_7656752519010 $T=48440 23850 0 0 $X=48360 $Y=23600
X16 67 M4_M3_CDNS_7656752519010 $T=53580 23850 0 0 $X=53500 $Y=23600
X17 53 M3_M2_CDNS_7656752519011 $T=150 23850 0 0 $X=70 $Y=23600
X18 54 M3_M2_CDNS_7656752519011 $T=5940 23850 0 0 $X=5860 $Y=23600
X19 5 M3_M2_CDNS_7656752519011 $T=9840 3330 0 0 $X=9760 $Y=3080
X20 55 M3_M2_CDNS_7656752519011 $T=16170 2650 0 0 $X=16090 $Y=2400
X21 56 M3_M2_CDNS_7656752519011 $T=16170 23850 0 0 $X=16090 $Y=23600
X22 57 M3_M2_CDNS_7656752519011 $T=21750 2650 0 0 $X=21670 $Y=2400
X23 58 M3_M2_CDNS_7656752519011 $T=21750 23850 0 0 $X=21670 $Y=23600
X24 59 M3_M2_CDNS_7656752519011 $T=26890 2650 0 0 $X=26810 $Y=2400
X25 60 M3_M2_CDNS_7656752519011 $T=26890 23850 0 0 $X=26810 $Y=23600
X26 61 M3_M2_CDNS_7656752519011 $T=32670 2650 0 0 $X=32590 $Y=2400
X27 62 M3_M2_CDNS_7656752519011 $T=32670 23850 0 0 $X=32590 $Y=23600
X28 63 M3_M2_CDNS_7656752519011 $T=40090 2650 0 0 $X=40010 $Y=2400
X29 64 M3_M2_CDNS_7656752519011 $T=40090 23850 0 0 $X=40010 $Y=23600
X30 65 M3_M2_CDNS_7656752519011 $T=48440 2650 0 0 $X=48360 $Y=2400
X31 66 M3_M2_CDNS_7656752519011 $T=48440 23850 0 0 $X=48360 $Y=23600
X32 67 M3_M2_CDNS_7656752519011 $T=53580 23850 0 0 $X=53500 $Y=23600
X33 2 M2_M1_CDNS_7656752519020 $T=4820 41440 0 0 $X=4740 $Y=41310
X34 10 M2_M1_CDNS_7656752519020 $T=13610 20240 0 0 $X=13530 $Y=20110
X35 11 M2_M1_CDNS_7656752519020 $T=13610 41440 0 0 $X=13530 $Y=41310
X36 16 M2_M1_CDNS_7656752519020 $T=19200 20240 0 0 $X=19120 $Y=20110
X37 17 M2_M1_CDNS_7656752519020 $T=19200 41440 0 0 $X=19120 $Y=41310
X38 23 M2_M1_CDNS_7656752519020 $T=31060 20240 0 0 $X=30980 $Y=20110
X39 22 M2_M1_CDNS_7656752519020 $T=31060 41440 0 0 $X=30980 $Y=41310
X40 24 M2_M1_CDNS_7656752519020 $T=31510 20240 0 0 $X=31430 $Y=20110
X41 25 M2_M1_CDNS_7656752519020 $T=31510 41440 0 0 $X=31430 $Y=41310
X42 34 M2_M1_CDNS_7656752519020 $T=40300 20240 0 0 $X=40220 $Y=20110
X43 35 M2_M1_CDNS_7656752519020 $T=40300 41440 0 0 $X=40220 $Y=41310
X44 36 M2_M1_CDNS_7656752519020 $T=45890 20240 0 0 $X=45810 $Y=20110
X45 37 M2_M1_CDNS_7656752519020 $T=45890 41440 0 0 $X=45810 $Y=41310
X46 45 M2_M1_CDNS_7656752519020 $T=57710 20240 0 0 $X=57630 $Y=20110
X47 46 M2_M1_CDNS_7656752519020 $T=57710 41440 0 0 $X=57630 $Y=41310
X48 52 M3_M2_CDNS_7656752519035 $T=560 24410 0 0 $X=480 $Y=24160
X49 68 M3_M2_CDNS_7656752519035 $T=9840 24410 0 0 $X=9760 $Y=24160
X50 69 M3_M2_CDNS_7656752519035 $T=17280 3210 0 0 $X=17200 $Y=2960
X51 70 M3_M2_CDNS_7656752519035 $T=17280 24410 0 0 $X=17200 $Y=24160
X52 71 M3_M2_CDNS_7656752519035 $T=22860 3210 0 0 $X=22780 $Y=2960
X53 72 M3_M2_CDNS_7656752519035 $T=22860 24410 0 0 $X=22780 $Y=24160
X54 73 M3_M2_CDNS_7656752519035 $T=27230 3210 0 0 $X=27150 $Y=2960
X55 74 M3_M2_CDNS_7656752519035 $T=27230 24410 0 0 $X=27150 $Y=24160
X56 75 M3_M2_CDNS_7656752519035 $T=36530 3210 0 0 $X=36450 $Y=2960
X57 76 M3_M2_CDNS_7656752519035 $T=36530 24410 0 0 $X=36450 $Y=24160
X58 77 M3_M2_CDNS_7656752519035 $T=43970 3210 0 0 $X=43890 $Y=2960
X59 78 M3_M2_CDNS_7656752519035 $T=43970 24410 0 0 $X=43890 $Y=24160
X60 79 M3_M2_CDNS_7656752519035 $T=49550 3210 0 0 $X=49470 $Y=2960
X61 80 M3_M2_CDNS_7656752519035 $T=49550 24410 0 0 $X=49470 $Y=24160
X62 52 M4_M3_CDNS_7656752519036 $T=560 24410 0 0 $X=480 $Y=24160
X63 5 M4_M3_CDNS_7656752519036 $T=9840 3330 0 0 $X=9760 $Y=3080
X64 68 M4_M3_CDNS_7656752519036 $T=9840 24410 0 0 $X=9760 $Y=24160
X65 69 M4_M3_CDNS_7656752519036 $T=17280 3210 0 0 $X=17200 $Y=2960
X66 70 M4_M3_CDNS_7656752519036 $T=17280 24410 0 0 $X=17200 $Y=24160
X67 71 M4_M3_CDNS_7656752519036 $T=22860 3210 0 0 $X=22780 $Y=2960
X68 72 M4_M3_CDNS_7656752519036 $T=22860 24410 0 0 $X=22780 $Y=24160
X69 73 M4_M3_CDNS_7656752519036 $T=27230 3210 0 0 $X=27150 $Y=2960
X70 74 M4_M3_CDNS_7656752519036 $T=27230 24410 0 0 $X=27150 $Y=24160
X71 75 M4_M3_CDNS_7656752519036 $T=36530 3210 0 0 $X=36450 $Y=2960
X72 76 M4_M3_CDNS_7656752519036 $T=36530 24410 0 0 $X=36450 $Y=24160
X73 77 M4_M3_CDNS_7656752519036 $T=43970 3210 0 0 $X=43890 $Y=2960
X74 78 M4_M3_CDNS_7656752519036 $T=43970 24410 0 0 $X=43890 $Y=24160
X75 79 M4_M3_CDNS_7656752519036 $T=49550 3210 0 0 $X=49470 $Y=2960
X76 80 M4_M3_CDNS_7656752519036 $T=49550 24410 0 0 $X=49470 $Y=24160
X77 53 M5_M4_CDNS_7656752519045 $T=150 23850 0 0 $X=70 $Y=23600
X78 54 M5_M4_CDNS_7656752519045 $T=5940 23850 0 0 $X=5860 $Y=23600
X79 55 M5_M4_CDNS_7656752519045 $T=16170 2650 0 0 $X=16090 $Y=2400
X80 56 M5_M4_CDNS_7656752519045 $T=16170 23850 0 0 $X=16090 $Y=23600
X81 57 M5_M4_CDNS_7656752519045 $T=21750 2650 0 0 $X=21670 $Y=2400
X82 58 M5_M4_CDNS_7656752519045 $T=21750 23850 0 0 $X=21670 $Y=23600
X83 59 M5_M4_CDNS_7656752519045 $T=26890 2650 0 0 $X=26810 $Y=2400
X84 60 M5_M4_CDNS_7656752519045 $T=26890 23850 0 0 $X=26810 $Y=23600
X85 61 M5_M4_CDNS_7656752519045 $T=32670 2650 0 0 $X=32590 $Y=2400
X86 62 M5_M4_CDNS_7656752519045 $T=32670 23850 0 0 $X=32590 $Y=23600
X87 63 M5_M4_CDNS_7656752519045 $T=40090 2650 0 0 $X=40010 $Y=2400
X88 64 M5_M4_CDNS_7656752519045 $T=40090 23850 0 0 $X=40010 $Y=23600
X89 65 M5_M4_CDNS_7656752519045 $T=48440 2650 0 0 $X=48360 $Y=2400
X90 66 M5_M4_CDNS_7656752519045 $T=48440 23850 0 0 $X=48360 $Y=23600
X91 67 M5_M4_CDNS_7656752519045 $T=53580 23850 0 0 $X=53500 $Y=23600
X92 53 M6_M5_CDNS_7656752519053 $T=150 23850 0 0 $X=70 $Y=23600
X93 54 M6_M5_CDNS_7656752519053 $T=5940 23850 0 0 $X=5860 $Y=23600
X94 55 M6_M5_CDNS_7656752519053 $T=16170 2650 0 0 $X=16090 $Y=2400
X95 56 M6_M5_CDNS_7656752519053 $T=16170 23850 0 0 $X=16090 $Y=23600
X96 57 M6_M5_CDNS_7656752519053 $T=21750 2650 0 0 $X=21670 $Y=2400
X97 58 M6_M5_CDNS_7656752519053 $T=21750 23850 0 0 $X=21670 $Y=23600
X98 59 M6_M5_CDNS_7656752519053 $T=26890 2650 0 0 $X=26810 $Y=2400
X99 60 M6_M5_CDNS_7656752519053 $T=26890 23850 0 0 $X=26810 $Y=23600
X100 61 M6_M5_CDNS_7656752519053 $T=32670 2650 0 0 $X=32590 $Y=2400
X101 62 M6_M5_CDNS_7656752519053 $T=32670 23850 0 0 $X=32590 $Y=23600
X102 63 M6_M5_CDNS_7656752519053 $T=40090 2650 0 0 $X=40010 $Y=2400
X103 64 M6_M5_CDNS_7656752519053 $T=40090 23850 0 0 $X=40010 $Y=23600
X104 65 M6_M5_CDNS_7656752519053 $T=48440 2650 0 0 $X=48360 $Y=2400
X105 66 M6_M5_CDNS_7656752519053 $T=48440 23850 0 0 $X=48360 $Y=23600
X106 67 M6_M5_CDNS_7656752519053 $T=53580 23850 0 0 $X=53500 $Y=23600
X107 81 M5_M4_CDNS_7656752519062 $T=9340 41110 0 0 $X=9120 $Y=40860
X108 82 M5_M4_CDNS_7656752519062 $T=18130 19910 0 0 $X=17910 $Y=19660
X109 83 M5_M4_CDNS_7656752519062 $T=18130 41110 0 0 $X=17910 $Y=40860
X110 84 M5_M4_CDNS_7656752519062 $T=23720 19910 0 0 $X=23500 $Y=19660
X111 85 M5_M4_CDNS_7656752519062 $T=23720 41110 0 0 $X=23500 $Y=40860
X112 86 M5_M4_CDNS_7656752519062 $T=26500 19910 0 0 $X=26280 $Y=19660
X113 87 M5_M4_CDNS_7656752519062 $T=26500 41110 0 0 $X=26280 $Y=40860
X114 88 M5_M4_CDNS_7656752519062 $T=36030 19910 0 0 $X=35810 $Y=19660
X115 89 M5_M4_CDNS_7656752519062 $T=36030 41110 0 0 $X=35810 $Y=40860
X116 90 M5_M4_CDNS_7656752519062 $T=44820 19910 0 0 $X=44600 $Y=19660
X117 91 M5_M4_CDNS_7656752519062 $T=44820 41110 0 0 $X=44600 $Y=40860
X118 92 M5_M4_CDNS_7656752519062 $T=50410 19910 0 0 $X=50190 $Y=19660
X119 93 M5_M4_CDNS_7656752519062 $T=50410 41110 0 0 $X=50190 $Y=40860
X120 94 M5_M4_CDNS_7656752519062 $T=53190 19910 0 0 $X=52970 $Y=19660
X121 95 M5_M4_CDNS_7656752519062 $T=53190 41110 0 0 $X=52970 $Y=40860
X122 81 M4_M3_CDNS_7656752519063 $T=9340 41110 0 0 $X=9120 $Y=40860
X123 82 M4_M3_CDNS_7656752519063 $T=18130 19910 0 0 $X=17910 $Y=19660
X124 83 M4_M3_CDNS_7656752519063 $T=18130 41110 0 0 $X=17910 $Y=40860
X125 84 M4_M3_CDNS_7656752519063 $T=23720 19910 0 0 $X=23500 $Y=19660
X126 85 M4_M3_CDNS_7656752519063 $T=23720 41110 0 0 $X=23500 $Y=40860
X127 86 M4_M3_CDNS_7656752519063 $T=26500 19910 0 0 $X=26280 $Y=19660
X128 87 M4_M3_CDNS_7656752519063 $T=26500 41110 0 0 $X=26280 $Y=40860
X129 88 M4_M3_CDNS_7656752519063 $T=36030 19910 0 0 $X=35810 $Y=19660
X130 89 M4_M3_CDNS_7656752519063 $T=36030 41110 0 0 $X=35810 $Y=40860
X131 90 M4_M3_CDNS_7656752519063 $T=44820 19910 0 0 $X=44600 $Y=19660
X132 91 M4_M3_CDNS_7656752519063 $T=44820 41110 0 0 $X=44600 $Y=40860
X133 92 M4_M3_CDNS_7656752519063 $T=50410 19910 0 0 $X=50190 $Y=19660
X134 93 M4_M3_CDNS_7656752519063 $T=50410 41110 0 0 $X=50190 $Y=40860
X135 94 M4_M3_CDNS_7656752519063 $T=53190 19910 0 0 $X=52970 $Y=19660
X136 95 M4_M3_CDNS_7656752519063 $T=53190 41110 0 0 $X=52970 $Y=40860
X137 81 M3_M2_CDNS_7656752519064 $T=9340 41110 0 0 $X=9120 $Y=40860
X138 82 M3_M2_CDNS_7656752519064 $T=18130 19910 0 0 $X=17910 $Y=19660
X139 83 M3_M2_CDNS_7656752519064 $T=18130 41110 0 0 $X=17910 $Y=40860
X140 84 M3_M2_CDNS_7656752519064 $T=23720 19910 0 0 $X=23500 $Y=19660
X141 85 M3_M2_CDNS_7656752519064 $T=23720 41110 0 0 $X=23500 $Y=40860
X142 86 M3_M2_CDNS_7656752519064 $T=26500 19910 0 0 $X=26280 $Y=19660
X143 87 M3_M2_CDNS_7656752519064 $T=26500 41110 0 0 $X=26280 $Y=40860
X144 88 M3_M2_CDNS_7656752519064 $T=36030 19910 0 0 $X=35810 $Y=19660
X145 89 M3_M2_CDNS_7656752519064 $T=36030 41110 0 0 $X=35810 $Y=40860
X146 90 M3_M2_CDNS_7656752519064 $T=44820 19910 0 0 $X=44600 $Y=19660
X147 91 M3_M2_CDNS_7656752519064 $T=44820 41110 0 0 $X=44600 $Y=40860
X148 92 M3_M2_CDNS_7656752519064 $T=50410 19910 0 0 $X=50190 $Y=19660
X149 93 M3_M2_CDNS_7656752519064 $T=50410 41110 0 0 $X=50190 $Y=40860
X150 94 M3_M2_CDNS_7656752519064 $T=53190 19910 0 0 $X=52970 $Y=19660
X151 95 M3_M2_CDNS_7656752519064 $T=53190 41110 0 0 $X=52970 $Y=40860
X152 81 M2_M1_CDNS_7656752519065 $T=9340 41110 0 0 $X=9120 $Y=40860
X153 82 M2_M1_CDNS_7656752519065 $T=18130 19910 0 0 $X=17910 $Y=19660
X154 83 M2_M1_CDNS_7656752519065 $T=18130 41110 0 0 $X=17910 $Y=40860
X155 84 M2_M1_CDNS_7656752519065 $T=23720 19910 0 0 $X=23500 $Y=19660
X156 85 M2_M1_CDNS_7656752519065 $T=23720 41110 0 0 $X=23500 $Y=40860
X157 86 M2_M1_CDNS_7656752519065 $T=26500 19910 0 0 $X=26280 $Y=19660
X158 87 M2_M1_CDNS_7656752519065 $T=26500 41110 0 0 $X=26280 $Y=40860
X159 88 M2_M1_CDNS_7656752519065 $T=36030 19910 0 0 $X=35810 $Y=19660
X160 89 M2_M1_CDNS_7656752519065 $T=36030 41110 0 0 $X=35810 $Y=40860
X161 90 M2_M1_CDNS_7656752519065 $T=44820 19910 0 0 $X=44600 $Y=19660
X162 91 M2_M1_CDNS_7656752519065 $T=44820 41110 0 0 $X=44600 $Y=40860
X163 92 M2_M1_CDNS_7656752519065 $T=50410 19910 0 0 $X=50190 $Y=19660
X164 93 M2_M1_CDNS_7656752519065 $T=50410 41110 0 0 $X=50190 $Y=40860
X165 94 M2_M1_CDNS_7656752519065 $T=53190 19910 0 0 $X=52970 $Y=19660
X166 95 M2_M1_CDNS_7656752519065 $T=53190 41110 0 0 $X=52970 $Y=40860
X167 81 M6_M5_CDNS_7656752519066 $T=9340 41110 0 0 $X=9120 $Y=40860
X168 82 M6_M5_CDNS_7656752519066 $T=18130 19910 0 0 $X=17910 $Y=19660
X169 83 M6_M5_CDNS_7656752519066 $T=18130 41110 0 0 $X=17910 $Y=40860
X170 84 M6_M5_CDNS_7656752519066 $T=23720 19910 0 0 $X=23500 $Y=19660
X171 85 M6_M5_CDNS_7656752519066 $T=23720 41110 0 0 $X=23500 $Y=40860
X172 86 M6_M5_CDNS_7656752519066 $T=26500 19910 0 0 $X=26280 $Y=19660
X173 87 M6_M5_CDNS_7656752519066 $T=26500 41110 0 0 $X=26280 $Y=40860
X174 88 M6_M5_CDNS_7656752519066 $T=36030 19910 0 0 $X=35810 $Y=19660
X175 89 M6_M5_CDNS_7656752519066 $T=36030 41110 0 0 $X=35810 $Y=40860
X176 90 M6_M5_CDNS_7656752519066 $T=44820 19910 0 0 $X=44600 $Y=19660
X177 91 M6_M5_CDNS_7656752519066 $T=44820 41110 0 0 $X=44600 $Y=40860
X178 92 M6_M5_CDNS_7656752519066 $T=50410 19910 0 0 $X=50190 $Y=19660
X179 93 M6_M5_CDNS_7656752519066 $T=50410 41110 0 0 $X=50190 $Y=40860
X180 94 M6_M5_CDNS_7656752519066 $T=53190 19910 0 0 $X=52970 $Y=19660
X181 95 M6_M5_CDNS_7656752519066 $T=53190 41110 0 0 $X=52970 $Y=40860
X182 7 2 4 3 81 110 186 AND $T=3670 43110 0 0 $X=4740 $Y=40010
X183 13 10 4 3 82 117 192 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X184 12 11 4 3 83 116 191 AND $T=12460 43110 0 0 $X=13530 $Y=40010
X185 21 16 4 3 84 123 198 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X186 20 17 4 3 85 122 197 AND $T=18050 43110 0 0 $X=19120 $Y=40010
X187 27 23 4 3 86 135 222 AND $T=32170 21910 1 180 $X=26920 $Y=18810
X188 26 22 4 3 87 134 221 AND $T=32170 43110 1 180 $X=26920 $Y=40010
X189 31 24 4 3 88 143 228 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X190 30 25 4 3 89 142 227 AND $T=30360 43110 0 0 $X=31430 $Y=40010
X191 39 34 4 3 90 149 236 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X192 38 35 4 3 91 148 235 AND $T=39150 43110 0 0 $X=40220 $Y=40010
X193 44 36 4 3 92 155 242 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X194 43 37 4 3 93 154 241 AND $T=44740 43110 0 0 $X=45810 $Y=40010
X195 48 45 4 3 94 162 249 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X196 47 46 4 3 95 161 248 AND $T=58860 43110 1 180 $X=53610 $Y=40010
X197 52 3 4 1 53 183 108 XOR $T=640 25900 1 0 $X=640 $Y=21200
X198 2 3 4 54 7 185 109 XOR $T=4740 40010 1 0 $X=4740 $Y=35310
X199 68 3 4 6 54 184 111 XOR $T=9740 25900 0 180 $X=6020 $Y=21200
X200 69 3 4 8 55 190 115 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X201 70 3 4 9 56 189 114 XOR $T=17180 25900 0 180 $X=13460 $Y=21200
X202 10 3 4 55 13 188 113 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X203 11 3 4 56 12 187 112 XOR $T=13530 40010 1 0 $X=13530 $Y=35310
X204 71 3 4 14 57 196 121 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X205 72 3 4 15 58 195 120 XOR $T=22760 25900 0 180 $X=19040 $Y=21200
X206 16 3 4 57 21 194 119 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X207 17 3 4 58 20 193 118 XOR $T=19120 40010 1 0 $X=19120 $Y=35310
X208 73 3 4 18 59 200 125 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X209 74 3 4 19 60 199 124 XOR $T=26810 25900 0 180 $X=23090 $Y=21200
X210 23 3 4 59 27 224 137 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X211 22 3 4 60 26 223 136 XOR $T=31140 40010 0 180 $X=27420 $Y=35310
X212 24 3 4 61 31 226 141 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X213 25 3 4 62 30 225 140 XOR $T=31430 40010 1 0 $X=31430 $Y=35310
X214 75 3 4 28 61 230 139 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X215 76 3 4 29 62 229 138 XOR $T=36470 25900 0 180 $X=32750 $Y=21200
X216 77 3 4 32 63 234 147 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X217 78 3 4 33 64 233 146 XOR $T=43890 25900 0 180 $X=40170 $Y=21200
X218 34 3 4 63 39 232 145 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X219 35 3 4 64 38 231 144 XOR $T=40220 40010 1 0 $X=40220 $Y=35310
X220 79 3 4 41 65 240 153 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X221 80 3 4 42 66 239 152 XOR $T=49450 25900 0 180 $X=45730 $Y=21200
X222 36 3 4 65 44 238 151 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X223 37 3 4 66 43 237 150 XOR $T=45810 40010 1 0 $X=45810 $Y=35310
X224 96 3 4 40 67 243 156 XOR $T=49650 25900 1 0 $X=49650 $Y=21200
X225 45 3 4 53 48 247 160 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X226 46 3 4 67 47 246 159 XOR $T=57790 40010 0 180 $X=54070 $Y=35310
X227 49 3 96 50 51 4 158 157 244 290
+ 291 245 HAdder $T=62720 27380 1 90 $X=53760 $Y=28180
X228 59 86 73 3 4 57 84 71 55 82
+ 69 97 5 98 99 104 105 106 107 260
+ 262 261 263 264 265 267 268 269 266 173
+ 174 177 178 176 179 180 175 181 182 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X229 60 87 74 3 4 58 85 72 56 83
+ 70 54 68 81 52 100 101 102 103 250
+ 252 251 253 254 255 257 258 259 256 163
+ 164 167 168 166 169 170 165 171 172 4bit_CLA_logic $T=26970 25900 1 180 $X=320 $Y=25900
X230 53 94 52 3 4 65 92 79 63 90
+ 77 61 75 88 73 130 131 132 133 280
+ 282 281 283 284 285 287 288 289 286 211
+ 212 215 216 214 217 218 213 219 220 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
X231 67 95 96 3 4 66 93 80 64 91
+ 78 62 76 89 74 126 127 128 129 270
+ 272 271 273 274 275 277 278 279 276 201
+ 202 205 206 204 207 208 203 209 210 4bit_CLA_logic $T=53660 25900 1 180 $X=27010 $Y=25900
M0 186 2 110 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5600 $Y=40350 $dt=0
M1 3 7 186 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5810 $Y=40350 $dt=0
M2 81 110 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=8230 $Y=40340 $dt=0
M3 192 10 117 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=19150 $dt=0
M4 191 11 116 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=40350 $dt=0
M5 3 13 192 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=19150 $dt=0
M6 3 12 191 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=40350 $dt=0
M7 82 117 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=19140 $dt=0
M8 83 116 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=40340 $dt=0
M9 198 16 123 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=19150 $dt=0
M10 197 17 122 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=40350 $dt=0
M11 3 21 198 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=19150 $dt=0
M12 3 20 197 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=40350 $dt=0
M13 84 123 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=19140 $dt=0
M14 85 122 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=40340 $dt=0
M15 3 135 86 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27520 $Y=19140 $dt=0
M16 3 134 87 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27520 $Y=40340 $dt=0
M17 222 27 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29940 $Y=19150 $dt=0
M18 221 26 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29940 $Y=40350 $dt=0
M19 135 23 222 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30150 $Y=19150 $dt=0
M20 134 22 221 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30150 $Y=40350 $dt=0
M21 228 24 143 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=19150 $dt=0
M22 227 25 142 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=40350 $dt=0
M23 3 31 228 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=19150 $dt=0
M24 3 30 227 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=40350 $dt=0
M25 88 143 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=19140 $dt=0
M26 89 142 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=40340 $dt=0
M27 236 34 149 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=19150 $dt=0
M28 235 35 148 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=40350 $dt=0
M29 3 39 236 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=19150 $dt=0
M30 3 38 235 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=40350 $dt=0
M31 90 149 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=19140 $dt=0
M32 91 148 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=40340 $dt=0
M33 242 36 155 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=19150 $dt=0
M34 241 37 154 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=40350 $dt=0
M35 3 44 242 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=19150 $dt=0
M36 3 43 241 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=40350 $dt=0
M37 92 155 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=19140 $dt=0
M38 93 154 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=40340 $dt=0
M39 3 162 94 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=19140 $dt=0
M40 3 161 95 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=40340 $dt=0
M41 249 48 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=19150 $dt=0
M42 248 47 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=40350 $dt=0
M43 162 45 249 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=19150 $dt=0
M44 161 46 248 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=40350 $dt=0
M45 4 107 99 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M46 4 103 52 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=34270 $dt=1
M47 183 52 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=22000 $dt=1
M48 266 98 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M49 256 81 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=34270 $dt=1
M50 1 53 52 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=22000 $dt=1
M51 183 108 1 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=22000 $dt=1
M52 4 53 108 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=22000 $dt=1
M53 185 2 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=36110 $dt=1
M54 110 2 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=5600 $Y=41790 $dt=1
M55 4 7 110 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=6010 $Y=41790 $dt=1
M56 54 7 2 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=36110 $dt=1
M57 111 54 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=22000 $dt=1
M58 185 109 54 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=36110 $dt=1
M59 6 111 184 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=22000 $dt=1
M60 4 7 109 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=36110 $dt=1
M61 81 110 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=8230 $Y=41600 $dt=1
M62 68 54 6 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=22000 $dt=1
M63 4 68 184 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=22000 $dt=1
M64 115 55 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M65 114 56 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=115.144 scb=0.0588049 scc=0.0138331 $X=13880 $Y=22000 $dt=1
M66 188 10 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M67 187 11 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=36110 $dt=1
M68 117 10 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.29 scb=0.029437 scc=0.00332952 $X=14390 $Y=20590 $dt=1
M69 116 11 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=14390 $Y=41790 $dt=1
M70 4 13 117 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=28.0435 scb=0.0261338 scc=0.00329543 $X=14800 $Y=20590 $dt=1
M71 4 12 116 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=14800 $Y=41790 $dt=1
M72 8 115 190 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M73 9 114 189 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.854 scb=0.0354545 scc=0.011187 $X=14810 $Y=22000 $dt=1
M74 55 13 10 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M75 56 12 11 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=36110 $dt=1
M76 69 55 8 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M77 70 56 9 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=15740 $Y=22000 $dt=1
M78 188 113 55 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M79 187 112 56 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=36110 $dt=1
M80 4 69 190 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M81 4 70 189 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=16670 $Y=22000 $dt=1
M82 4 13 113 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M83 4 12 112 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=36110 $dt=1
M84 82 117 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=17020 $Y=20400 $dt=1
M85 83 116 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=17020 $Y=41600 $dt=1
M86 121 57 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M87 120 58 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=19460 $Y=22000 $dt=1
M88 194 16 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M89 193 17 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=36110 $dt=1
M90 123 16 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=19980 $Y=20590 $dt=1
M91 122 17 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=19980 $Y=41790 $dt=1
M92 14 121 196 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M93 4 21 123 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=20390 $Y=20590 $dt=1
M94 15 120 195 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=20390 $Y=22000 $dt=1
M95 4 20 122 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=20390 $Y=41790 $dt=1
M96 57 21 16 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M97 58 20 17 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=36110 $dt=1
M98 71 57 14 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M99 72 58 15 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=21320 $Y=22000 $dt=1
M100 194 119 57 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M101 193 118 58 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=36110 $dt=1
M102 4 71 196 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M103 4 72 195 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=22250 $Y=22000 $dt=1
M104 4 21 119 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M105 4 20 118 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=36110 $dt=1
M106 84 123 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=22610 $Y=20400 $dt=1
M107 85 122 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=22610 $Y=41600 $dt=1
M108 125 59 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M109 124 60 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=23510 $Y=22000 $dt=1
M110 18 125 200 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M111 19 124 199 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=24440 $Y=22000 $dt=1
M112 73 59 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M113 74 60 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=25370 $Y=22000 $dt=1
M114 4 73 200 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M115 4 74 199 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=26300 $Y=22000 $dt=1
M116 4 133 73 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M117 4 129 74 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=34270 $dt=1
M118 4 135 86 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=27520 $Y=20400 $dt=1
M119 4 134 87 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=27520 $Y=41600 $dt=1
M120 137 27 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M121 136 26 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=36110 $dt=1
M122 286 88 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M123 276 89 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=34270 $dt=1
M124 59 137 224 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M125 60 136 223 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=36110 $dt=1
M126 23 27 59 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M127 22 26 60 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=36110 $dt=1
M128 135 27 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=29740 $Y=20590 $dt=1
M129 134 26 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=29740 $Y=41790 $dt=1
M130 4 23 135 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=30150 $Y=20590 $dt=1
M131 4 22 134 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=30150 $Y=41790 $dt=1
M132 4 23 224 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M133 4 22 223 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=36110 $dt=1
M134 226 24 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M135 225 25 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=36110 $dt=1
M136 143 24 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32290 $Y=20590 $dt=1
M137 142 25 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=32290 $Y=41790 $dt=1
M138 4 31 143 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32700 $Y=20590 $dt=1
M139 4 30 142 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=32700 $Y=41790 $dt=1
M140 61 31 24 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M141 62 30 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=36110 $dt=1
M142 139 61 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M143 138 62 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=33170 $Y=22000 $dt=1
M144 226 141 61 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M145 225 140 62 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=36110 $dt=1
M146 28 139 230 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M147 29 138 229 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=34100 $Y=22000 $dt=1
M148 4 31 141 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M149 4 30 140 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=36110 $dt=1
M150 88 143 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=34920 $Y=20400 $dt=1
M151 89 142 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=34920 $Y=41600 $dt=1
M152 75 61 28 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M153 76 62 29 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35030 $Y=22000 $dt=1
M154 4 75 230 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M155 4 76 229 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35960 $Y=22000 $dt=1
M156 147 63 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M157 146 64 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=40590 $Y=22000 $dt=1
M158 232 34 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M159 231 35 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=36110 $dt=1
M160 149 34 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41080 $Y=20590 $dt=1
M161 148 35 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=41080 $Y=41790 $dt=1
M162 4 39 149 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41490 $Y=20590 $dt=1
M163 4 38 148 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=41490 $Y=41790 $dt=1
M164 32 147 234 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M165 33 146 233 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=41520 $Y=22000 $dt=1
M166 63 39 34 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M167 64 38 35 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=36110 $dt=1
M168 77 63 32 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M169 78 64 33 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=42450 $Y=22000 $dt=1
M170 232 145 63 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M171 231 144 64 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=36110 $dt=1
M172 4 77 234 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M173 4 78 233 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=43380 $Y=22000 $dt=1
M174 4 39 145 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M175 4 38 144 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=36110 $dt=1
M176 90 149 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=43710 $Y=20400 $dt=1
M177 91 148 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=43710 $Y=41600 $dt=1
M178 153 65 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M179 152 66 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=46150 $Y=22000 $dt=1
M180 238 36 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M181 237 37 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=36110 $dt=1
M182 155 36 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=46670 $Y=20590 $dt=1
M183 154 37 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=46670 $Y=41790 $dt=1
M184 41 153 240 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M185 4 44 155 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=47080 $Y=20590 $dt=1
M186 42 152 239 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=47080 $Y=22000 $dt=1
M187 4 43 154 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.816 scb=0.0254064 scc=0.0032946 $X=47080 $Y=41790 $dt=1
M188 65 44 36 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M189 66 43 37 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=36110 $dt=1
M190 79 65 41 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=48010 $Y=800 $dt=1
M191 80 66 42 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48010 $Y=22000 $dt=1
M192 238 151 65 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M193 237 150 66 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=36110 $dt=1
M194 4 79 240 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=48940 $Y=800 $dt=1
M195 4 80 239 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48940 $Y=22000 $dt=1
M196 4 44 151 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M197 4 43 150 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=36110 $dt=1
M198 92 155 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=49300 $Y=20400 $dt=1
M199 93 154 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=49300 $Y=41600 $dt=1
M200 243 96 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=50070 $Y=22000 $dt=1
M201 40 67 96 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51000 $Y=22000 $dt=1
M202 243 156 40 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51930 $Y=22000 $dt=1
M203 4 67 156 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=52860 $Y=22000 $dt=1
M204 4 162 94 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=54210 $Y=20400 $dt=1
M205 4 161 95 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8162 scb=0.0285373 scc=0.00672168 $X=54210 $Y=41600 $dt=1
M206 160 48 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M207 159 47 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=36110 $dt=1
M208 53 160 247 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M209 67 159 246 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=36110 $dt=1
M210 291 158 96 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=55830 $Y=32900 $dt=1
M211 4 157 291 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56040 $Y=32900 $dt=1
M212 45 48 53 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M213 46 47 67 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=36110 $dt=1
M214 162 48 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=29.0043 scb=0.0273456 scc=0.00330147 $X=56430 $Y=20590 $dt=1
M215 161 47 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=28.969 scb=0.0273266 scc=0.00330146 $X=56430 $Y=41790 $dt=1
M216 4 45 162 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=33.5338 scb=0.0350848 scc=0.00355838 $X=56840 $Y=20590 $dt=1
M217 4 46 161 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=33.4985 scb=0.0350659 scc=0.00355836 $X=56840 $Y=41790 $dt=1
M218 4 157 290 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56970 $Y=32900 $dt=1
M219 4 45 247 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M220 4 46 246 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=36110 $dt=1
M221 290 158 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57380 $Y=32900 $dt=1
M222 49 51 290 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57790 $Y=32900 $dt=1
M223 290 50 49 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=58200 $Y=32900 $dt=1
M224 4 50 157 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=59130 $Y=32900 $dt=1
M225 4 51 158 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=60060 $Y=32900 $dt=1
.ends MAC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceProjectMAC                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceProjectMAC 199 198 197 196 195 194 193 192 191 200
+ 201 202 203 204 205 206 239 235 230 226
+ 222 220 214 236 234 229 225 221 219 213
+ 210 237 47 238 232 227 223 217 215 211
+ 208 231 233 228 224 218 216 212 209 207
+ 147 116 67 141 115 87 133 131 144 65
+ 140 78 76 77 66 117 83
** N=838 EP=67 FDC=2230
X0 1 M5_M4_CDNS_765675251900 $T=8680 96730 0 0 $X=8600 $Y=96600
X1 2 M5_M4_CDNS_765675251900 $T=17180 99960 0 0 $X=17100 $Y=99830
X2 3 M5_M4_CDNS_765675251900 $T=21730 98530 0 0 $X=21650 $Y=98400
X3 4 M5_M4_CDNS_765675251900 $T=25170 119910 0 0 $X=25090 $Y=119780
X4 5 M5_M4_CDNS_765675251900 $T=41900 93630 0 0 $X=41820 $Y=93500
X5 6 M5_M4_CDNS_765675251900 $T=42370 94030 0 0 $X=42290 $Y=93900
X6 7 M5_M4_CDNS_765675251900 $T=43570 92930 0 0 $X=43490 $Y=92800
X7 8 M5_M4_CDNS_765675251900 $T=43920 95730 0 0 $X=43840 $Y=95600
X8 9 M5_M4_CDNS_765675251900 $T=45720 98250 0 0 $X=45640 $Y=98120
X9 1 M5_M4_CDNS_765675251901 $T=8680 95430 0 0 $X=8550 $Y=95300
X10 10 M5_M4_CDNS_765675251901 $T=16520 72380 0 0 $X=16390 $Y=72250
X11 11 M5_M4_CDNS_765675251901 $T=19630 96730 0 0 $X=19500 $Y=96600
X12 8 M5_M4_CDNS_765675251901 $T=43920 101770 0 0 $X=43790 $Y=101640
X13 12 M4_M3_CDNS_765675251902 $T=2330 93930 0 0 $X=2200 $Y=93850
X14 13 M4_M3_CDNS_765675251902 $T=2680 98180 0 0 $X=2550 $Y=98100
X15 14 M4_M3_CDNS_765675251902 $T=6790 81230 0 0 $X=6660 $Y=81150
X16 15 M4_M3_CDNS_765675251902 $T=7630 101030 0 0 $X=7500 $Y=100950
X17 16 M4_M3_CDNS_765675251902 $T=8330 95080 0 0 $X=8200 $Y=95000
X18 1 M4_M3_CDNS_765675251902 $T=8680 95430 0 0 $X=8550 $Y=95350
X19 17 M4_M3_CDNS_765675251902 $T=9030 96030 0 0 $X=8900 $Y=95950
X20 8 M4_M3_CDNS_765675251902 $T=9730 95730 0 0 $X=9600 $Y=95650
X21 18 M4_M3_CDNS_765675251902 $T=10080 94280 0 0 $X=9950 $Y=94200
X22 7 M4_M3_CDNS_765675251902 $T=12540 92930 0 0 $X=12410 $Y=92850
X23 19 M4_M3_CDNS_765675251902 $T=15020 98900 0 0 $X=14890 $Y=98820
X24 5 M4_M3_CDNS_765675251902 $T=15890 93630 0 0 $X=15760 $Y=93550
X25 10 M4_M3_CDNS_765675251902 $T=16520 72380 0 0 $X=16390 $Y=72300
X26 20 M4_M3_CDNS_765675251902 $T=16890 86180 0 0 $X=16760 $Y=86100
X27 21 M4_M3_CDNS_765675251902 $T=17310 93230 0 0 $X=17180 $Y=93150
X28 12 M4_M3_CDNS_765675251902 $T=17310 93930 0 0 $X=17180 $Y=93850
X29 18 M4_M3_CDNS_765675251902 $T=17310 94280 0 0 $X=17180 $Y=94200
X30 22 M4_M3_CDNS_765675251902 $T=17310 94630 0 0 $X=17180 $Y=94550
X31 17 M4_M3_CDNS_765675251902 $T=17310 96030 0 0 $X=17180 $Y=95950
X32 23 M4_M3_CDNS_765675251902 $T=18510 99620 0 0 $X=18380 $Y=99540
X33 2 M4_M3_CDNS_765675251902 $T=18670 88620 0 0 $X=18540 $Y=88540
X34 24 M4_M3_CDNS_765675251902 $T=18930 99580 0 0 $X=18800 $Y=99500
X35 6 M4_M3_CDNS_765675251902 $T=19890 98480 0 0 $X=19760 $Y=98400
X36 23 M4_M3_CDNS_765675251902 $T=20680 81120 0 0 $X=20550 $Y=81040
X37 3 M4_M3_CDNS_765675251902 $T=22430 98530 0 0 $X=22300 $Y=98450
X38 25 M4_M3_CDNS_765675251902 $T=24660 97130 0 0 $X=24530 $Y=97050
X39 26 M4_M3_CDNS_765675251902 $T=25200 109890 0 0 $X=25070 $Y=109810
X40 27 M4_M3_CDNS_765675251902 $T=25740 97130 0 0 $X=25610 $Y=97050
X41 28 M4_M3_CDNS_765675251902 $T=25910 97830 0 0 $X=25780 $Y=97750
X42 29 M4_M3_CDNS_765675251902 $T=26000 113050 0 0 $X=25870 $Y=112970
X43 30 M4_M3_CDNS_765675251902 $T=27040 100570 0 0 $X=26910 $Y=100490
X44 31 M4_M3_CDNS_765675251902 $T=27410 101330 0 0 $X=27280 $Y=101250
X45 13 M4_M3_CDNS_765675251902 $T=29840 98180 0 0 $X=29710 $Y=98100
X46 19 M4_M3_CDNS_765675251902 $T=30510 93230 0 0 $X=30380 $Y=93150
X47 15 M4_M3_CDNS_765675251902 $T=31330 101030 0 0 $X=31200 $Y=100950
X48 32 M4_M3_CDNS_765675251902 $T=34650 79520 0 0 $X=34520 $Y=79440
X49 32 M4_M3_CDNS_765675251902 $T=34650 101010 0 0 $X=34520 $Y=100930
X50 33 M4_M3_CDNS_765675251902 $T=35310 99930 0 0 $X=35180 $Y=99850
X51 20 M4_M3_CDNS_765675251902 $T=37310 86180 0 0 $X=37180 $Y=86100
X52 34 M4_M3_CDNS_765675251902 $T=39310 85830 0 0 $X=39180 $Y=85750
X53 35 M4_M3_CDNS_765675251902 $T=40690 94330 0 0 $X=40560 $Y=94250
X54 11 M4_M3_CDNS_765675251902 $T=41190 96030 0 0 $X=41060 $Y=95950
X55 36 M4_M3_CDNS_765675251902 $T=42140 100630 0 0 $X=42010 $Y=100550
X56 24 M4_M3_CDNS_765675251902 $T=46090 99580 0 0 $X=45960 $Y=99500
X57 37 M4_M3_CDNS_765675251902 $T=46480 100160 0 0 $X=46350 $Y=100080
X58 38 M4_M3_CDNS_765675251902 $T=48490 98880 0 0 $X=48360 $Y=98800
X59 19 M5_M4_CDNS_765675251903 $T=15020 98900 0 0 $X=14890 $Y=98530
X60 10 M5_M4_CDNS_765675251903 $T=16520 91390 0 0 $X=16390 $Y=91020
X61 39 M5_M4_CDNS_765675251903 $T=16830 118300 0 0 $X=16700 $Y=117930
X62 40 M5_M4_CDNS_765675251903 $T=17570 117850 0 0 $X=17440 $Y=117480
X63 2 M5_M4_CDNS_765675251903 $T=18670 88620 0 0 $X=18540 $Y=88250
X64 40 M5_M4_CDNS_765675251903 $T=21030 80000 0 0 $X=20900 $Y=79630
X65 4 M5_M4_CDNS_765675251903 $T=25170 72590 0 0 $X=25040 $Y=72220
X66 32 M5_M4_CDNS_765675251903 $T=34650 79520 0 0 $X=34520 $Y=79150
X67 5 M5_M4_CDNS_765675251903 $T=41900 100280 0 0 $X=41770 $Y=99910
X68 6 M5_M4_CDNS_765675251903 $T=42370 100280 0 0 $X=42240 $Y=99910
X69 7 M5_M4_CDNS_765675251903 $T=43570 102040 0 0 $X=43440 $Y=101670
X70 21 M4_M3_CDNS_765675251904 $T=1900 93230 0 0 $X=1820 $Y=93100
X71 41 M4_M3_CDNS_765675251904 $T=3650 92530 0 0 $X=3570 $Y=92400
X72 42 M4_M3_CDNS_765675251904 $T=5880 82250 0 0 $X=5800 $Y=82120
X73 42 M4_M3_CDNS_765675251904 $T=5880 87300 0 0 $X=5800 $Y=87170
X74 43 M4_M3_CDNS_765675251904 $T=8380 96380 0 0 $X=8300 $Y=96250
X75 30 M4_M3_CDNS_765675251904 $T=10800 100570 0 0 $X=10720 $Y=100440
X76 44 M4_M3_CDNS_765675251904 $T=11190 74080 0 0 $X=11110 $Y=73950
X77 10 M4_M3_CDNS_765675251904 $T=16520 91390 0 0 $X=16440 $Y=91260
X78 2 M4_M3_CDNS_765675251904 $T=17180 100220 0 0 $X=17100 $Y=100090
X79 39 M4_M3_CDNS_765675251904 $T=21380 73000 0 0 $X=21300 $Y=72870
X80 45 M4_M3_CDNS_765675251904 $T=31390 100680 0 0 $X=31310 $Y=100550
X81 41 M4_M3_CDNS_765675251904 $T=41800 92530 0 0 $X=41720 $Y=92400
X82 9 M4_M3_CDNS_765675251904 $T=45720 98510 0 0 $X=45640 $Y=98380
X83 46 M4_M3_CDNS_765675251904 $T=47260 97130 0 0 $X=47180 $Y=97000
X84 31 M4_M3_CDNS_765675251904 $T=55100 101330 0 0 $X=55020 $Y=101200
X85 47 M4_M3_CDNS_765675251904 $T=59240 48070 0 90 $X=59110 $Y=47990
X86 28 M4_M3_CDNS_765675251904 $T=59910 100550 0 0 $X=59830 $Y=100420
X87 22 M4_M3_CDNS_765675251905 $T=-390 94630 0 0 $X=-520 $Y=94260
X88 9 M4_M3_CDNS_765675251905 $T=3030 97480 0 0 $X=2900 $Y=97110
X89 48 M4_M3_CDNS_765675251905 $T=8310 71930 0 0 $X=8180 $Y=71560
X90 44 M4_M3_CDNS_765675251905 $T=11190 88980 0 0 $X=11060 $Y=88610
X91 29 M4_M3_CDNS_765675251905 $T=13830 111740 0 0 $X=13700 $Y=111370
X92 39 M4_M3_CDNS_765675251905 $T=16830 118300 0 0 $X=16700 $Y=117930
X93 38 M4_M3_CDNS_765675251905 $T=17310 98880 0 0 $X=17180 $Y=98510
X94 40 M4_M3_CDNS_765675251905 $T=17570 117850 0 0 $X=17440 $Y=117480
X95 33 M4_M3_CDNS_765675251905 $T=17580 99930 0 0 $X=17450 $Y=99560
X96 49 M4_M3_CDNS_765675251905 $T=18930 101770 0 0 $X=18800 $Y=101400
X97 35 M4_M3_CDNS_765675251905 $T=20130 103160 0 0 $X=20000 $Y=102790
X98 3 M4_M3_CDNS_765675251905 $T=20130 111380 0 0 $X=20000 $Y=111010
X99 50 M4_M3_CDNS_765675251905 $T=22690 99230 0 0 $X=22560 $Y=98860
X100 4 M4_M3_CDNS_765675251905 $T=25170 72590 0 0 $X=25040 $Y=72220
X101 43 M4_M3_CDNS_765675251905 $T=41190 100330 0 0 $X=41060 $Y=99960
X102 5 M4_M3_CDNS_765675251905 $T=41900 100280 0 0 $X=41770 $Y=99910
X103 6 M4_M3_CDNS_765675251905 $T=42370 100280 0 0 $X=42240 $Y=99910
X104 16 M4_M3_CDNS_765675251905 $T=42400 95080 0 0 $X=42270 $Y=94710
X105 37 M4_M3_CDNS_765675251905 $T=43230 100160 0 0 $X=43100 $Y=99790
X106 7 M4_M3_CDNS_765675251905 $T=43570 102040 0 0 $X=43440 $Y=101670
X107 34 M4_M3_CDNS_765675251905 $T=47850 88280 0 0 $X=47720 $Y=87910
X108 51 M3_M2_CDNS_765675251906 $T=1330 80160 0 0 $X=1250 $Y=80030
X109 51 M3_M2_CDNS_765675251906 $T=1330 104390 0 0 $X=1250 $Y=104260
X110 26 M3_M2_CDNS_765675251906 $T=2250 111070 0 0 $X=2170 $Y=110940
X111 26 M3_M2_CDNS_765675251906 $T=2250 112040 0 0 $X=2170 $Y=111910
X112 13 M3_M2_CDNS_765675251906 $T=2680 88600 0 0 $X=2600 $Y=88470
X113 9 M3_M2_CDNS_765675251906 $T=3030 97480 0 0 $X=2950 $Y=97350
X114 45 M3_M2_CDNS_765675251906 $T=4510 82980 0 0 $X=4430 $Y=82850
X115 52 M3_M2_CDNS_765675251906 $T=5010 87930 0 0 $X=4930 $Y=87800
X116 15 M3_M2_CDNS_765675251906 $T=6280 95080 0 0 $X=6200 $Y=94950
X117 16 M3_M2_CDNS_765675251906 $T=8330 95660 0 0 $X=8250 $Y=95530
X118 17 M3_M2_CDNS_765675251906 $T=9030 100590 0 0 $X=8950 $Y=100460
X119 8 M3_M2_CDNS_765675251906 $T=9730 98040 0 0 $X=9650 $Y=97910
X120 44 M3_M2_CDNS_765675251906 $T=11190 88980 0 0 $X=11110 $Y=88850
X121 53 M3_M2_CDNS_765675251906 $T=11410 96380 0 0 $X=11330 $Y=96250
X122 54 M3_M2_CDNS_765675251906 $T=11710 95430 0 0 $X=11630 $Y=95300
X123 54 M3_M2_CDNS_765675251906 $T=11710 97340 0 0 $X=11630 $Y=97210
X124 54 M3_M2_CDNS_765675251906 $T=11710 99520 0 0 $X=11630 $Y=99390
X125 7 M3_M2_CDNS_765675251906 $T=12540 94390 0 0 $X=12460 $Y=94260
X126 5 M3_M2_CDNS_765675251906 $T=15890 94270 0 0 $X=15810 $Y=94140
X127 39 M3_M2_CDNS_765675251906 $T=16830 118300 0 0 $X=16750 $Y=118170
X128 55 M3_M2_CDNS_765675251906 $T=16920 74000 0 0 $X=16840 $Y=73870
X129 1 M3_M2_CDNS_765675251906 $T=17100 96730 0 0 $X=17020 $Y=96600
X130 40 M3_M2_CDNS_765675251906 $T=17570 117850 0 0 $X=17490 $Y=117720
X131 33 M3_M2_CDNS_765675251906 $T=17580 99930 0 0 $X=17500 $Y=99800
X132 49 M3_M2_CDNS_765675251906 $T=18140 98310 0 0 $X=18060 $Y=98180
X133 49 M3_M2_CDNS_765675251906 $T=18140 99650 0 0 $X=18060 $Y=99520
X134 56 M3_M2_CDNS_765675251906 $T=21690 86530 0 0 $X=21610 $Y=86400
X135 34 M3_M2_CDNS_765675251906 $T=22040 85830 0 0 $X=21960 $Y=85700
X136 3 M3_M2_CDNS_765675251906 $T=22430 96730 0 0 $X=22350 $Y=96600
X137 50 M3_M2_CDNS_765675251906 $T=22690 99230 0 0 $X=22610 $Y=99100
X138 30 M3_M2_CDNS_765675251906 $T=27040 100380 0 0 $X=26960 $Y=100250
X139 31 M3_M2_CDNS_765675251906 $T=27410 98880 0 0 $X=27330 $Y=98750
X140 1 M3_M2_CDNS_765675251906 $T=29350 98980 0 0 $X=29270 $Y=98850
X141 19 M3_M2_CDNS_765675251906 $T=30510 93570 0 0 $X=30430 $Y=93440
X142 57 M3_M2_CDNS_765675251906 $T=31450 90030 0 0 $X=31370 $Y=89900
X143 42 M3_M2_CDNS_765675251906 $T=32290 87300 0 0 $X=32210 $Y=87170
X144 58 M3_M2_CDNS_765675251906 $T=35660 72840 0 0 $X=35580 $Y=72710
X145 59 M3_M2_CDNS_765675251906 $T=36230 101110 0 0 $X=36150 $Y=100980
X146 59 M3_M2_CDNS_765675251906 $T=36230 104400 0 0 $X=36150 $Y=104270
X147 60 M3_M2_CDNS_765675251906 $T=38790 101400 0 0 $X=38710 $Y=101270
X148 17 M3_M2_CDNS_765675251906 $T=39890 96030 0 0 $X=39810 $Y=95900
X149 35 M3_M2_CDNS_765675251906 $T=40690 96080 0 0 $X=40610 $Y=95950
X150 41 M3_M2_CDNS_765675251906 $T=41800 96430 0 0 $X=41720 $Y=96300
X151 16 M3_M2_CDNS_765675251906 $T=42400 95250 0 0 $X=42320 $Y=95120
X152 7 M3_M2_CDNS_765675251906 $T=43570 102040 0 0 $X=43490 $Y=101910
X153 8 M3_M2_CDNS_765675251906 $T=43920 101770 0 0 $X=43840 $Y=101640
X154 24 M3_M2_CDNS_765675251906 $T=46090 100580 0 0 $X=46010 $Y=100450
X155 61 M3_M2_CDNS_765675251906 $T=46110 91130 0 0 $X=46030 $Y=91000
X156 37 M3_M2_CDNS_765675251906 $T=46480 98530 0 0 $X=46400 $Y=98400
X157 62 M3_M2_CDNS_765675251906 $T=47390 96330 0 0 $X=47310 $Y=96200
X158 34 M3_M2_CDNS_765675251906 $T=47850 88280 0 0 $X=47770 $Y=88150
X159 38 M3_M2_CDNS_765675251906 $T=48490 99650 0 0 $X=48410 $Y=99520
X160 27 M3_M2_CDNS_765675251906 $T=49320 97160 0 0 $X=49240 $Y=97030
X161 31 M3_M2_CDNS_765675251906 $T=55100 100540 0 0 $X=55020 $Y=100410
X162 28 M3_M2_CDNS_765675251906 $T=59910 100810 0 0 $X=59830 $Y=100680
X163 37 M3_M2_CDNS_765675251906 $T=60410 97860 0 0 $X=60330 $Y=97730
X164 63 M3_M2_CDNS_765675251906 $T=60710 100630 0 0 $X=60630 $Y=100500
X165 19 M5_M4_CDNS_765675251907 $T=17730 94630 0 0 $X=17600 $Y=94550
X166 6 M5_M4_CDNS_765675251907 $T=19280 94030 0 0 $X=19150 $Y=93950
X167 6 M5_M4_CDNS_765675251907 $T=19280 98480 0 0 $X=19150 $Y=98400
X168 11 M5_M4_CDNS_765675251907 $T=19630 96030 0 0 $X=19500 $Y=95950
X169 23 M5_M4_CDNS_765675251907 $T=19980 81120 0 0 $X=19850 $Y=81040
X170 39 M5_M4_CDNS_765675251907 $T=21380 89430 0 0 $X=21250 $Y=89350
X171 3 M5_M4_CDNS_765675251907 $T=21730 111380 0 0 $X=21600 $Y=111300
X172 25 M5_M4_CDNS_765675251907 $T=24660 90430 0 0 $X=24530 $Y=90350
X173 19 M5_M4_CDNS_765675251907 $T=30510 94630 0 0 $X=30380 $Y=94550
X174 45 M5_M4_CDNS_765675251907 $T=31390 100230 0 0 $X=31260 $Y=100150
X175 36 M5_M4_CDNS_765675251907 $T=33310 100630 0 0 $X=33180 $Y=100550
X176 35 M5_M4_CDNS_765675251907 $T=40690 103160 0 0 $X=40560 $Y=103080
X177 43 M5_M4_CDNS_765675251907 $T=41190 96380 0 0 $X=41060 $Y=96300
X178 9 M5_M4_CDNS_765675251907 $T=45720 97480 0 0 $X=45590 $Y=97400
X179 64 M5_M4_CDNS_765675251908 $T=18230 111270 0 0 $X=18150 $Y=111020
X180 64 M5_M4_CDNS_765675251908 $T=20330 89330 0 0 $X=20250 $Y=89080
X181 2 M2_M1_CDNS_765675251909 $T=17180 111020 0 0 $X=17100 $Y=110770
X182 64 M2_M1_CDNS_765675251909 $T=18230 111270 0 0 $X=18150 $Y=111020
X183 49 M2_M1_CDNS_765675251909 $T=37450 101760 0 0 $X=37370 $Y=101510
X184 65 M2_M1_CDNS_765675251909 $T=40310 37330 0 0 $X=40230 $Y=37080
X185 47 M2_M1_CDNS_765675251909 $T=60710 26810 0 0 $X=60630 $Y=26560
X186 66 M4_M3_CDNS_7656752519010 $T=4820 42750 0 0 $X=4740 $Y=42500
X187 64 M4_M3_CDNS_7656752519010 $T=18230 111270 0 0 $X=18150 $Y=111020
X188 65 M4_M3_CDNS_7656752519010 $T=40310 37330 0 0 $X=40230 $Y=37080
X189 67 M4_M3_CDNS_7656752519010 $T=60960 21490 0 0 $X=60880 $Y=21240
X190 65 M4_M3_CDNS_7656752519010 $T=61270 38260 0 0 $X=61190 $Y=38010
X191 2 M3_M2_CDNS_7656752519011 $T=17180 111020 0 0 $X=17100 $Y=110770
X192 64 M3_M2_CDNS_7656752519011 $T=18230 111270 0 0 $X=18150 $Y=111020
X193 49 M3_M2_CDNS_7656752519011 $T=37450 101760 0 0 $X=37370 $Y=101510
X194 65 M3_M2_CDNS_7656752519011 $T=40310 37330 0 0 $X=40230 $Y=37080
X195 47 M3_M2_CDNS_7656752519011 $T=60710 26810 0 0 $X=60630 $Y=26560
X196 23 M5_M4_CDNS_7656752519012 $T=18510 99620 0 0 $X=18140 $Y=99490
X197 50 M5_M4_CDNS_7656752519012 $T=22690 99230 0 0 $X=22320 $Y=99100
X198 25 M5_M4_CDNS_7656752519012 $T=24660 97130 0 0 $X=24290 $Y=97000
X199 19 M5_M4_CDNS_7656752519012 $T=30510 93230 0 0 $X=30140 $Y=93100
X200 32 M5_M4_CDNS_7656752519012 $T=34650 101010 0 0 $X=34280 $Y=100880
X201 35 M5_M4_CDNS_7656752519012 $T=40690 94330 0 0 $X=40320 $Y=94200
X202 43 M5_M4_CDNS_7656752519012 $T=41190 100330 0 0 $X=40820 $Y=100200
X203 20 M4_M3_CDNS_7656752519013 $T=16890 88280 0 0 $X=16760 $Y=88150
X204 1 M4_M3_CDNS_7656752519013 $T=17100 96730 0 0 $X=16970 $Y=96600
X205 11 M4_M3_CDNS_7656752519013 $T=19630 96730 0 0 $X=19500 $Y=96600
X206 40 M4_M3_CDNS_7656752519013 $T=21030 80000 0 0 $X=20900 $Y=79870
X207 46 M4_M3_CDNS_7656752519013 $T=21270 96780 0 0 $X=21140 $Y=96650
X208 8 M4_M3_CDNS_7656752519013 $T=43920 101770 0 0 $X=43790 $Y=101640
X209 68 M3_M2_CDNS_7656752519014 $T=-700 73550 0 0 $X=-830 $Y=73180
X210 22 M3_M2_CDNS_7656752519014 $T=-390 94630 0 0 $X=-520 $Y=94260
X211 69 M3_M2_CDNS_7656752519014 $T=3160 89330 0 0 $X=3030 $Y=88960
X212 41 M3_M2_CDNS_7656752519014 $T=3650 90320 0 0 $X=3520 $Y=89950
X213 36 M3_M2_CDNS_7656752519014 $T=4000 89680 0 0 $X=3870 $Y=89310
X214 42 M3_M2_CDNS_7656752519014 $T=5880 81840 0 0 $X=5750 $Y=81470
X215 14 M3_M2_CDNS_7656752519014 $T=6580 110930 0 0 $X=6450 $Y=110560
X216 1 M3_M2_CDNS_7656752519014 $T=8790 112270 0 0 $X=8660 $Y=111900
X217 32 M3_M2_CDNS_7656752519014 $T=9930 79520 0 0 $X=9800 $Y=79150
X218 25 M3_M2_CDNS_7656752519014 $T=9950 90030 0 0 $X=9820 $Y=89660
X219 18 M3_M2_CDNS_7656752519014 $T=9950 111680 0 0 $X=9820 $Y=111310
X220 30 M3_M2_CDNS_7656752519014 $T=10800 97220 0 0 $X=10670 $Y=96850
X221 29 M3_M2_CDNS_7656752519014 $T=13830 111740 0 0 $X=13700 $Y=111370
X222 19 M3_M2_CDNS_7656752519014 $T=15160 111350 0 0 $X=15030 $Y=110980
X223 23 M3_M2_CDNS_7656752519014 $T=17880 118160 0 0 $X=17750 $Y=117790
X224 49 M3_M2_CDNS_7656752519014 $T=18930 101770 0 0 $X=18800 $Y=101400
X225 11 M3_M2_CDNS_7656752519014 $T=19630 96730 0 0 $X=19500 $Y=96360
X226 6 M3_M2_CDNS_7656752519014 $T=20550 98480 0 0 $X=20420 $Y=98110
X227 46 M3_M2_CDNS_7656752519014 $T=21270 96780 0 0 $X=21140 $Y=96410
X228 2 M3_M2_CDNS_7656752519014 $T=21290 88620 0 0 $X=21160 $Y=88250
X229 26 M3_M2_CDNS_7656752519014 $T=25200 101440 0 0 $X=25070 $Y=101070
X230 52 M3_M2_CDNS_7656752519014 $T=25520 88380 0 0 $X=25390 $Y=88010
X231 29 M3_M2_CDNS_7656752519014 $T=26000 101440 0 0 $X=25870 $Y=101070
X232 70 M3_M2_CDNS_7656752519014 $T=31890 98160 0 0 $X=31760 $Y=97790
X233 71 M3_M2_CDNS_7656752519014 $T=32630 79950 0 0 $X=32500 $Y=79580
X234 32 M3_M2_CDNS_7656752519014 $T=34650 101460 0 0 $X=34520 $Y=101090
X235 13 M3_M2_CDNS_7656752519014 $T=36630 99550 0 0 $X=36500 $Y=99180
X236 57 M3_M2_CDNS_7656752519014 $T=36860 88380 0 0 $X=36730 $Y=88010
X237 63 M3_M2_CDNS_7656752519014 $T=36940 96980 0 0 $X=36810 $Y=96610
X238 72 M3_M2_CDNS_7656752519014 $T=39070 97510 0 0 $X=38940 $Y=97140
X239 37 M3_M2_CDNS_7656752519014 $T=43230 100160 0 0 $X=43100 $Y=99790
X240 56 M3_M2_CDNS_7656752519014 $T=47850 80600 0 0 $X=47720 $Y=80230
X241 62 M3_M2_CDNS_7656752519014 $T=55310 88680 0 0 $X=55180 $Y=88310
X242 70 M3_M2_CDNS_7656752519014 $T=57720 100570 0 0 $X=57590 $Y=100200
X243 21 M3_M2_CDNS_7656752519017 $T=1900 111430 0 0 $X=1770 $Y=111350
X244 50 M3_M2_CDNS_7656752519017 $T=2490 82630 0 0 $X=2360 $Y=82550
X245 14 M3_M2_CDNS_7656752519017 $T=6580 95430 0 0 $X=6450 $Y=95350
X246 14 M3_M2_CDNS_7656752519017 $T=6790 89980 0 0 $X=6660 $Y=89900
X247 44 M3_M2_CDNS_7656752519017 $T=7280 95430 0 0 $X=7150 $Y=95350
X248 44 M3_M2_CDNS_7656752519017 $T=7280 107040 0 0 $X=7150 $Y=106960
X249 48 M3_M2_CDNS_7656752519017 $T=8310 71930 0 0 $X=8180 $Y=71850
X250 73 M3_M2_CDNS_7656752519017 $T=8960 90460 0 0 $X=8830 $Y=90380
X251 44 M3_M2_CDNS_7656752519017 $T=11190 71410 0 0 $X=11060 $Y=71330
X252 74 M3_M2_CDNS_7656752519017 $T=12880 91070 0 0 $X=12750 $Y=90990
X253 69 M3_M2_CDNS_7656752519017 $T=13310 89330 0 0 $X=13180 $Y=89250
X254 58 M3_M2_CDNS_7656752519017 $T=16450 81790 0 0 $X=16320 $Y=81710
X255 1 M3_M2_CDNS_7656752519017 $T=17100 95130 0 0 $X=16970 $Y=95050
X256 38 M3_M2_CDNS_7656752519017 $T=17310 98880 0 0 $X=17180 $Y=98800
X257 75 M3_M2_CDNS_7656752519017 $T=18260 80900 0 0 $X=18130 $Y=80820
X258 24 M3_M2_CDNS_7656752519017 $T=18930 99230 0 0 $X=18800 $Y=99150
X259 76 M3_M2_CDNS_7656752519017 $T=19250 38020 0 0 $X=19120 $Y=37940
X260 75 M3_M2_CDNS_7656752519017 $T=19940 80900 0 0 $X=19810 $Y=80820
X261 58 M3_M2_CDNS_7656752519017 $T=20310 81790 0 0 $X=20180 $Y=81710
X262 61 M3_M2_CDNS_7656752519017 $T=20540 91130 0 0 $X=20410 $Y=91050
X263 71 M3_M2_CDNS_7656752519017 $T=20680 80600 0 0 $X=20550 $Y=80520
X264 40 M3_M2_CDNS_7656752519017 $T=21030 80000 0 0 $X=20900 $Y=79920
X265 3 M3_M2_CDNS_7656752519017 $T=22430 95730 0 0 $X=22300 $Y=95650
X266 10 M3_M2_CDNS_7656752519017 $T=23880 90830 0 0 $X=23750 $Y=90750
X267 18 M3_M2_CDNS_7656752519017 $T=24330 94280 0 0 $X=24200 $Y=94200
X268 27 M3_M2_CDNS_7656752519017 $T=25170 97130 0 0 $X=25040 $Y=97050
X269 25 M3_M2_CDNS_7656752519017 $T=27010 96830 0 0 $X=26880 $Y=96750
X270 48 M3_M2_CDNS_7656752519017 $T=28680 91830 0 0 $X=28550 $Y=91750
X271 1 M3_M2_CDNS_7656752519017 $T=29350 95130 0 0 $X=29220 $Y=95050
X272 1 M3_M2_CDNS_7656752519017 $T=29350 101440 0 0 $X=29220 $Y=101360
X273 21 M3_M2_CDNS_7656752519017 $T=29800 93230 0 0 $X=29670 $Y=93150
X274 3 M3_M2_CDNS_7656752519017 $T=31030 95730 0 0 $X=30900 $Y=95650
X275 45 M3_M2_CDNS_7656752519017 $T=31170 100680 0 0 $X=31040 $Y=100600
X276 15 M3_M2_CDNS_7656752519017 $T=31610 101030 0 0 $X=31480 $Y=100950
X277 71 M3_M2_CDNS_7656752519017 $T=32630 80600 0 0 $X=32500 $Y=80520
X278 12 M3_M2_CDNS_7656752519017 $T=33720 93930 0 0 $X=33590 $Y=93850
X279 54 M3_M2_CDNS_7656752519017 $T=35430 95430 0 0 $X=35300 $Y=95350
X280 58 M3_M2_CDNS_7656752519017 $T=35660 81440 0 0 $X=35530 $Y=81360
X281 53 M3_M2_CDNS_7656752519017 $T=35830 96380 0 0 $X=35700 $Y=96300
X282 73 M3_M2_CDNS_7656752519017 $T=36510 90460 0 0 $X=36380 $Y=90380
X283 20 M3_M2_CDNS_7656752519017 $T=37310 88780 0 0 $X=37180 $Y=88700
X284 22 M3_M2_CDNS_7656752519017 $T=39490 94630 0 0 $X=39360 $Y=94550
X285 33 M3_M2_CDNS_7656752519017 $T=40290 99930 0 0 $X=40160 $Y=99850
X286 43 M3_M2_CDNS_7656752519017 $T=41190 100330 0 0 $X=41060 $Y=100250
X287 11 M3_M2_CDNS_7656752519017 $T=41450 96030 0 0 $X=41320 $Y=95950
X288 5 M3_M2_CDNS_7656752519017 $T=41900 100280 0 0 $X=41770 $Y=100200
X289 36 M3_M2_CDNS_7656752519017 $T=42400 100630 0 0 $X=42270 $Y=100550
X290 37 M3_M2_CDNS_7656752519017 $T=46480 97860 0 0 $X=46350 $Y=97780
X291 46 M3_M2_CDNS_7656752519017 $T=46830 97130 0 0 $X=46700 $Y=97050
X292 72 M3_M2_CDNS_7656752519017 $T=52950 97510 0 0 $X=52820 $Y=97430
X293 77 M5_M4_CDNS_7656752519018 $T=13070 42750 0 0 $X=12820 $Y=42670
X294 50 M5_M4_CDNS_7656752519018 $T=22690 82630 0 0 $X=22440 $Y=82550
X295 36 M5_M4_CDNS_7656752519018 $T=29310 89680 0 0 $X=29060 $Y=89600
X296 45 M5_M4_CDNS_7656752519018 $T=31390 82980 0 0 $X=31140 $Y=82900
X297 26 M4_M3_CDNS_7656752519019 $T=230 110810 0 0 $X=-20 $Y=110730
X298 76 M4_M3_CDNS_7656752519019 $T=18650 42750 0 0 $X=18400 $Y=42670
X299 50 M4_M3_CDNS_7656752519019 $T=22690 82630 0 0 $X=22440 $Y=82550
X300 48 M4_M3_CDNS_7656752519019 $T=28680 91830 0 0 $X=28430 $Y=91750
X301 36 M4_M3_CDNS_7656752519019 $T=29310 89680 0 0 $X=29060 $Y=89600
X302 45 M4_M3_CDNS_7656752519019 $T=31390 82980 0 0 $X=31140 $Y=82900
X303 78 M4_M3_CDNS_7656752519019 $T=54600 47040 0 0 $X=54350 $Y=46960
X304 68 M2_M1_CDNS_7656752519020 $T=-700 118270 0 0 $X=-780 $Y=118140
X305 79 M2_M1_CDNS_7656752519020 $T=-80 103430 0 0 $X=-160 $Y=103300
X306 68 M2_M1_CDNS_7656752519020 $T=1280 120900 0 0 $X=1200 $Y=120770
X307 13 M2_M1_CDNS_7656752519020 $T=1560 88600 0 0 $X=1480 $Y=88470
X308 26 M2_M1_CDNS_7656752519020 $T=2130 112300 0 0 $X=2050 $Y=112170
X309 50 M2_M1_CDNS_7656752519020 $T=2490 80510 0 0 $X=2410 $Y=80380
X310 9 M2_M1_CDNS_7656752519020 $T=2510 97480 0 0 $X=2430 $Y=97350
X311 80 M2_M1_CDNS_7656752519020 $T=2550 97970 0 0 $X=2470 $Y=97840
X312 52 M2_M1_CDNS_7656752519020 $T=2830 91250 0 0 $X=2750 $Y=91120
X313 79 M2_M1_CDNS_7656752519020 $T=2870 103430 0 0 $X=2790 $Y=103300
X314 81 M2_M1_CDNS_7656752519020 $T=3160 104950 0 0 $X=3080 $Y=104820
X315 82 M2_M1_CDNS_7656752519020 $T=3210 73020 0 0 $X=3130 $Y=72890
X316 83 M2_M1_CDNS_7656752519020 $T=3240 120790 0 0 $X=3160 $Y=120660
X317 81 M2_M1_CDNS_7656752519020 $T=3540 110950 0 0 $X=3460 $Y=110820
X318 41 M2_M1_CDNS_7656752519020 $T=3650 90320 0 0 $X=3570 $Y=90190
X319 45 M2_M1_CDNS_7656752519020 $T=4510 82170 0 0 $X=4430 $Y=82040
X320 71 M2_M1_CDNS_7656752519020 $T=5550 73490 0 0 $X=5470 $Y=73360
X321 83 M2_M1_CDNS_7656752519020 $T=6150 121230 0 0 $X=6070 $Y=121100
X322 84 M2_M1_CDNS_7656752519020 $T=6540 96610 0 0 $X=6460 $Y=96480
X323 84 M2_M1_CDNS_7656752519020 $T=6540 105070 0 0 $X=6460 $Y=104940
X324 14 M2_M1_CDNS_7656752519020 $T=6580 110930 0 0 $X=6500 $Y=110800
X325 75 M2_M1_CDNS_7656752519020 $T=6890 80900 0 0 $X=6810 $Y=80770
X326 16 M2_M1_CDNS_7656752519020 $T=8330 96510 0 0 $X=8250 $Y=96380
X327 43 M2_M1_CDNS_7656752519020 $T=8380 97010 0 0 $X=8300 $Y=96880
X328 71 M2_M1_CDNS_7656752519020 $T=8420 79410 0 0 $X=8340 $Y=79280
X329 1 M2_M1_CDNS_7656752519020 $T=8790 112270 0 0 $X=8710 $Y=112140
X330 47 M2_M1_CDNS_7656752519020 $T=8900 120860 0 0 $X=8820 $Y=120730
X331 8 M2_M1_CDNS_7656752519020 $T=9210 98040 0 0 $X=9130 $Y=97910
X332 25 M2_M1_CDNS_7656752519020 $T=9950 90030 0 0 $X=9870 $Y=89900
X333 18 M2_M1_CDNS_7656752519020 $T=9950 111680 0 0 $X=9870 $Y=111550
X334 44 M2_M1_CDNS_7656752519020 $T=10550 120910 0 0 $X=10470 $Y=120780
X335 53 M2_M1_CDNS_7656752519020 $T=11410 97340 0 0 $X=11330 $Y=97210
X336 53 M2_M1_CDNS_7656752519020 $T=11410 104450 0 0 $X=11330 $Y=104320
X337 47 M2_M1_CDNS_7656752519020 $T=11820 121150 0 0 $X=11740 $Y=121020
X338 7 M2_M1_CDNS_7656752519020 $T=12540 96660 0 0 $X=12460 $Y=96530
X339 74 M2_M1_CDNS_7656752519020 $T=12880 82460 0 0 $X=12800 $Y=82330
X340 39 M2_M1_CDNS_7656752519020 $T=13220 120920 0 0 $X=13140 $Y=120790
X341 44 M2_M1_CDNS_7656752519020 $T=13830 71410 0 0 $X=13750 $Y=71280
X342 29 M2_M1_CDNS_7656752519020 $T=13830 111740 0 0 $X=13750 $Y=111610
X343 83 M2_M1_CDNS_7656752519020 $T=14580 120890 0 0 $X=14500 $Y=120760
X344 83 M2_M1_CDNS_7656752519020 $T=15410 120950 0 0 $X=15330 $Y=120820
X345 85 M2_M1_CDNS_7656752519020 $T=15840 90790 0 0 $X=15760 $Y=90660
X346 5 M2_M1_CDNS_7656752519020 $T=15890 96510 0 0 $X=15810 $Y=96380
X347 40 M2_M1_CDNS_7656752519020 $T=16200 120910 0 0 $X=16120 $Y=120780
X348 86 M2_M1_CDNS_7656752519020 $T=16370 79450 0 0 $X=16290 $Y=79320
X349 86 M2_M1_CDNS_7656752519020 $T=17860 71590 0 0 $X=17780 $Y=71460
X350 86 M2_M1_CDNS_7656752519020 $T=17860 75760 0 0 $X=17780 $Y=75630
X351 23 M2_M1_CDNS_7656752519020 $T=18910 120910 0 0 $X=18830 $Y=120780
X352 87 M2_M1_CDNS_7656752519020 $T=19440 17190 0 0 $X=19360 $Y=17060
X353 11 M2_M1_CDNS_7656752519020 $T=19630 96660 0 0 $X=19550 $Y=96530
X354 3 M2_M1_CDNS_7656752519020 $T=20130 111380 0 0 $X=20050 $Y=111250
X355 47 M2_M1_CDNS_7656752519020 $T=20250 120910 0 0 $X=20170 $Y=120780
X356 61 M2_M1_CDNS_7656752519020 $T=20540 90800 0 0 $X=20460 $Y=90670
X357 6 M2_M1_CDNS_7656752519020 $T=20550 98480 0 0 $X=20470 $Y=98350
X358 56 M2_M1_CDNS_7656752519020 $T=20620 91480 0 0 $X=20540 $Y=91350
X359 46 M2_M1_CDNS_7656752519020 $T=21270 96660 0 0 $X=21190 $Y=96530
X360 2 M2_M1_CDNS_7656752519020 $T=21290 88620 0 0 $X=21210 $Y=88490
X361 39 M2_M1_CDNS_7656752519020 $T=21380 72640 0 0 $X=21300 $Y=72510
X362 4 M2_M1_CDNS_7656752519020 $T=21890 120910 0 0 $X=21810 $Y=120780
X363 34 M2_M1_CDNS_7656752519020 $T=22040 88140 0 0 $X=21960 $Y=88010
X364 88 M2_M1_CDNS_7656752519020 $T=22380 111680 0 0 $X=22300 $Y=111550
X365 59 M2_M1_CDNS_7656752519020 $T=22680 104400 0 0 $X=22600 $Y=104270
X366 47 M2_M1_CDNS_7656752519020 $T=23170 121220 0 0 $X=23090 $Y=121090
X367 10 M2_M1_CDNS_7656752519020 $T=23880 96990 0 0 $X=23800 $Y=96860
X368 18 M2_M1_CDNS_7656752519020 $T=24330 96980 0 0 $X=24250 $Y=96850
X369 4 M2_M1_CDNS_7656752519020 $T=25170 72590 0 0 $X=25090 $Y=72460
X370 26 M2_M1_CDNS_7656752519020 $T=25200 101440 0 0 $X=25120 $Y=101310
X371 52 M2_M1_CDNS_7656752519020 $T=25520 88380 0 0 $X=25440 $Y=88250
X372 89 M2_M1_CDNS_7656752519020 $T=25910 81790 0 0 $X=25830 $Y=81660
X373 29 M2_M1_CDNS_7656752519020 $T=26000 101440 0 0 $X=25920 $Y=101310
X374 31 M2_M1_CDNS_7656752519020 $T=26330 98880 0 0 $X=26250 $Y=98750
X375 88 M2_M1_CDNS_7656752519020 $T=26400 101440 0 0 $X=26320 $Y=101310
X376 50 M2_M1_CDNS_7656752519020 $T=26660 100640 0 0 $X=26580 $Y=100510
X377 25 M2_M1_CDNS_7656752519020 $T=27220 96830 0 0 $X=27140 $Y=96700
X378 85 M2_M1_CDNS_7656752519020 $T=27600 97880 0 0 $X=27520 $Y=97750
X379 48 M2_M1_CDNS_7656752519020 $T=28680 99330 0 0 $X=28600 $Y=99200
X380 21 M2_M1_CDNS_7656752519020 $T=29800 99700 0 0 $X=29720 $Y=99570
X381 90 M2_M1_CDNS_7656752519020 $T=30580 79400 0 0 $X=30500 $Y=79270
X382 3 M2_M1_CDNS_7656752519020 $T=31030 99380 0 0 $X=30950 $Y=99250
X383 91 M2_M1_CDNS_7656752519020 $T=31470 98510 0 0 $X=31390 $Y=98380
X384 15 M2_M1_CDNS_7656752519020 $T=31820 101030 0 0 $X=31740 $Y=100900
X385 92 M2_M1_CDNS_7656752519020 $T=31890 89330 0 0 $X=31810 $Y=89200
X386 42 M2_M1_CDNS_7656752519020 $T=32290 88570 0 0 $X=32210 $Y=88440
X387 71 M2_M1_CDNS_7656752519020 $T=32630 79950 0 0 $X=32550 $Y=79820
X388 12 M2_M1_CDNS_7656752519020 $T=33720 96520 0 0 $X=33640 $Y=96390
X389 58 M2_M1_CDNS_7656752519020 $T=35660 72580 0 0 $X=35580 $Y=72450
X390 59 M2_M1_CDNS_7656752519020 $T=36230 100850 0 0 $X=36150 $Y=100720
X391 73 M2_M1_CDNS_7656752519020 $T=36510 90170 0 0 $X=36430 $Y=90040
X392 13 M2_M1_CDNS_7656752519020 $T=36630 99550 0 0 $X=36550 $Y=99420
X393 57 M2_M1_CDNS_7656752519020 $T=36860 88380 0 0 $X=36780 $Y=88250
X394 63 M2_M1_CDNS_7656752519020 $T=36940 96980 0 0 $X=36860 $Y=96850
X395 30 M2_M1_CDNS_7656752519020 $T=37020 100380 0 0 $X=36940 $Y=100250
X396 60 M2_M1_CDNS_7656752519020 $T=38790 100280 0 0 $X=38710 $Y=100150
X397 72 M2_M1_CDNS_7656752519020 $T=39070 97510 0 0 $X=38990 $Y=97380
X398 22 M2_M1_CDNS_7656752519020 $T=39490 97070 0 0 $X=39410 $Y=96940
X399 93 M2_M1_CDNS_7656752519020 $T=39570 89330 0 0 $X=39490 $Y=89200
X400 17 M2_M1_CDNS_7656752519020 $T=39890 96740 0 0 $X=39810 $Y=96610
X401 33 M2_M1_CDNS_7656752519020 $T=40290 100140 0 0 $X=40210 $Y=100010
X402 35 M2_M1_CDNS_7656752519020 $T=40690 96700 0 0 $X=40610 $Y=96570
X403 94 M2_M1_CDNS_7656752519020 $T=40910 81680 0 0 $X=40830 $Y=81550
X404 95 M2_M1_CDNS_7656752519020 $T=40910 90200 0 0 $X=40830 $Y=90070
X405 41 M2_M1_CDNS_7656752519020 $T=41090 98880 0 0 $X=41010 $Y=98750
X406 43 M2_M1_CDNS_7656752519020 $T=41490 100330 0 0 $X=41410 $Y=100200
X407 5 M2_M1_CDNS_7656752519020 $T=41900 100920 0 0 $X=41820 $Y=100790
X408 11 M2_M1_CDNS_7656752519020 $T=42280 101440 0 0 $X=42200 $Y=101310
X409 6 M2_M1_CDNS_7656752519020 $T=42370 100280 0 0 $X=42290 $Y=100150
X410 96 M2_M1_CDNS_7656752519020 $T=43230 81310 0 0 $X=43150 $Y=81180
X411 37 M2_M1_CDNS_7656752519020 $T=43230 100160 0 0 $X=43150 $Y=100030
X412 97 M2_M1_CDNS_7656752519020 $T=43250 63930 0 0 $X=43170 $Y=63800
X413 7 M2_M1_CDNS_7656752519020 $T=43570 101180 0 0 $X=43490 $Y=101050
X414 20 M2_M1_CDNS_7656752519020 $T=43970 88780 0 0 $X=43890 $Y=88650
X415 98 M2_M1_CDNS_7656752519020 $T=43970 97220 0 0 $X=43890 $Y=97090
X416 36 M2_M1_CDNS_7656752519020 $T=45790 100630 0 0 $X=45710 $Y=100500
X417 24 M2_M1_CDNS_7656752519020 $T=46570 101430 0 0 $X=46490 $Y=101300
X418 46 M2_M1_CDNS_7656752519020 $T=46830 100430 0 0 $X=46750 $Y=100300
X419 62 M2_M1_CDNS_7656752519020 $T=47390 100770 0 0 $X=47310 $Y=100640
X420 99 M2_M1_CDNS_7656752519020 $T=47850 97220 0 0 $X=47770 $Y=97090
X421 100 M2_M1_CDNS_7656752519020 $T=47870 72330 0 0 $X=47790 $Y=72200
X422 101 M2_M1_CDNS_7656752519020 $T=48520 63930 0 0 $X=48440 $Y=63800
X423 94 M2_M1_CDNS_7656752519020 $T=48590 81680 0 0 $X=48510 $Y=81550
X424 102 M2_M1_CDNS_7656752519020 $T=48600 97620 0 0 $X=48520 $Y=97490
X425 103 M2_M1_CDNS_7656752519020 $T=50910 71610 0 0 $X=50830 $Y=71480
X426 104 M2_M1_CDNS_7656752519020 $T=50910 82090 0 0 $X=50830 $Y=81960
X427 105 M2_M1_CDNS_7656752519020 $T=50910 88980 0 0 $X=50830 $Y=88850
X428 106 M2_M1_CDNS_7656752519020 $T=50910 100060 0 0 $X=50830 $Y=99930
X429 60 M2_M1_CDNS_7656752519020 $T=51300 101460 0 0 $X=51220 $Y=101330
X430 98 M2_M1_CDNS_7656752519020 $T=51700 99890 0 0 $X=51620 $Y=99760
X431 99 M2_M1_CDNS_7656752519020 $T=52090 101040 0 0 $X=52010 $Y=100910
X432 107 M2_M1_CDNS_7656752519020 $T=54160 79510 0 0 $X=54080 $Y=79380
X433 107 M2_M1_CDNS_7656752519020 $T=54160 81970 0 0 $X=54080 $Y=81840
X434 9 M2_M1_CDNS_7656752519020 $T=54300 101520 0 0 $X=54220 $Y=101390
X435 108 M2_M1_CDNS_7656752519020 $T=54500 97910 0 0 $X=54420 $Y=97780
X436 105 M2_M1_CDNS_7656752519020 $T=54570 88980 0 0 $X=54490 $Y=88850
X437 31 M2_M1_CDNS_7656752519020 $T=55100 100280 0 0 $X=55020 $Y=100150
X438 62 M2_M1_CDNS_7656752519020 $T=55310 88680 0 0 $X=55230 $Y=88550
X439 72 M2_M1_CDNS_7656752519020 $T=55910 99800 0 0 $X=55830 $Y=99670
X440 108 M2_M1_CDNS_7656752519020 $T=56300 100030 0 0 $X=56220 $Y=99900
X441 109 M2_M1_CDNS_7656752519020 $T=56420 80850 0 0 $X=56340 $Y=80720
X442 110 M2_M1_CDNS_7656752519020 $T=56700 100940 0 0 $X=56620 $Y=100810
X443 111 M2_M1_CDNS_7656752519020 $T=57090 99720 0 0 $X=57010 $Y=99590
X444 112 M2_M1_CDNS_7656752519020 $T=59200 71290 0 0 $X=59120 $Y=71160
X445 113 M2_M1_CDNS_7656752519020 $T=59200 98490 0 0 $X=59120 $Y=98360
X446 114 M2_M1_CDNS_7656752519020 $T=59210 88110 0 0 $X=59130 $Y=87980
X447 28 M2_M1_CDNS_7656752519020 $T=59910 101100 0 0 $X=59830 $Y=100970
X448 63 M2_M1_CDNS_7656752519020 $T=60710 100970 0 0 $X=60630 $Y=100840
X449 37 M2_M1_CDNS_7656752519020 $T=61110 100660 0 0 $X=61030 $Y=100530
X450 115 M3_M2_CDNS_7656752519021 $T=7600 46120 0 0 $X=7230 $Y=45990
X451 43 M3_M2_CDNS_7656752519021 $T=8380 97010 0 0 $X=8010 $Y=96880
X452 10 M3_M2_CDNS_7656752519021 $T=16310 72380 0 0 $X=15940 $Y=72250
X453 20 M3_M2_CDNS_7656752519021 $T=16890 88280 0 0 $X=16520 $Y=88150
X454 67 M3_M2_CDNS_7656752519021 $T=20370 44250 0 0 $X=20000 $Y=44120
X455 55 M3_M2_CDNS_7656752519021 $T=20550 72330 0 0 $X=20180 $Y=72200
X456 116 M3_M2_CDNS_7656752519021 $T=24280 44200 0 0 $X=23910 $Y=44070
X457 4 M3_M2_CDNS_7656752519021 $T=25170 72590 0 0 $X=24800 $Y=72460
X458 23 M3_M2_CDNS_7656752519021 $T=25170 80000 0 0 $X=24800 $Y=79870
X459 117 M3_M2_CDNS_7656752519021 $T=34080 44250 0 0 $X=33710 $Y=44120
X460 68 M2_M1_CDNS_7656752519023 $T=-700 73550 0 0 $X=-830 $Y=73470
X461 22 M2_M1_CDNS_7656752519023 $T=-390 94630 0 0 $X=-520 $Y=94550
X462 22 M2_M1_CDNS_7656752519023 $T=-390 111110 0 0 $X=-520 $Y=111030
X463 79 M2_M1_CDNS_7656752519023 $T=-80 65150 0 0 $X=-210 $Y=65070
X464 118 M2_M1_CDNS_7656752519023 $T=230 71260 0 0 $X=100 $Y=71180
X465 22 M2_M1_CDNS_7656752519023 $T=1380 111110 0 0 $X=1250 $Y=111030
X466 48 M2_M1_CDNS_7656752519023 $T=2510 71930 0 0 $X=2380 $Y=71850
X467 51 M2_M1_CDNS_7656752519023 $T=2550 104900 0 0 $X=2420 $Y=104820
X468 21 M2_M1_CDNS_7656752519023 $T=2620 111430 0 0 $X=2490 $Y=111350
X469 79 M2_M1_CDNS_7656752519023 $T=3160 65150 0 0 $X=3030 $Y=65070
X470 69 M2_M1_CDNS_7656752519023 $T=3160 89330 0 0 $X=3030 $Y=89250
X471 36 M2_M1_CDNS_7656752519023 $T=4000 89680 0 0 $X=3870 $Y=89600
X472 10 M2_M1_CDNS_7656752519023 $T=4110 72380 0 0 $X=3980 $Y=72300
X473 38 M2_M1_CDNS_7656752519023 $T=4200 96710 0 0 $X=4070 $Y=96630
X474 42 M2_M1_CDNS_7656752519023 $T=5880 81840 0 0 $X=5750 $Y=81760
X475 119 M2_M1_CDNS_7656752519023 $T=5910 103750 0 0 $X=5780 $Y=103670
X476 118 M2_M1_CDNS_7656752519023 $T=6530 71260 0 0 $X=6400 $Y=71180
X477 84 M2_M1_CDNS_7656752519023 $T=6540 82200 0 0 $X=6410 $Y=82120
X478 73 M2_M1_CDNS_7656752519023 $T=7650 90460 0 0 $X=7520 $Y=90380
X479 71 M2_M1_CDNS_7656752519023 $T=8420 80300 0 0 $X=8290 $Y=80220
X480 15 M2_M1_CDNS_7656752519023 $T=8790 89080 0 0 $X=8660 $Y=89000
X481 17 M2_M1_CDNS_7656752519023 $T=8790 100590 0 0 $X=8660 $Y=100510
X482 58 M2_M1_CDNS_7656752519023 $T=9230 81790 0 0 $X=9100 $Y=81710
X483 68 M2_M1_CDNS_7656752519023 $T=9710 73550 0 0 $X=9580 $Y=73470
X484 32 M2_M1_CDNS_7656752519023 $T=9930 79520 0 0 $X=9800 $Y=79440
X485 54 M2_M1_CDNS_7656752519023 $T=9950 99520 0 0 $X=9820 $Y=99440
X486 120 M2_M1_CDNS_7656752519023 $T=10020 72080 0 0 $X=9890 $Y=72000
X487 30 M2_M1_CDNS_7656752519023 $T=10800 97220 0 0 $X=10670 $Y=97140
X488 53 M2_M1_CDNS_7656752519023 $T=13830 104450 0 0 $X=13700 $Y=104370
X489 51 M2_M1_CDNS_7656752519023 $T=13850 79870 0 0 $X=13720 $Y=79790
X490 55 M2_M1_CDNS_7656752519023 $T=13890 74000 0 0 $X=13760 $Y=73920
X491 121 M2_M1_CDNS_7656752519023 $T=13890 82600 0 0 $X=13760 $Y=82520
X492 120 M2_M1_CDNS_7656752519023 $T=14570 72080 0 0 $X=14440 $Y=72000
X493 24 M2_M1_CDNS_7656752519023 $T=14570 99230 0 0 $X=14440 $Y=99150
X494 33 M2_M1_CDNS_7656752519023 $T=14990 99930 0 0 $X=14860 $Y=99850
X495 19 M2_M1_CDNS_7656752519023 $T=15160 111350 0 0 $X=15030 $Y=111270
X496 49 M2_M1_CDNS_7656752519023 $T=15540 97390 0 0 $X=15410 $Y=97310
X497 20 M2_M1_CDNS_7656752519023 $T=16890 88280 0 0 $X=16760 $Y=88200
X498 122 M2_M1_CDNS_7656752519023 $T=18230 72030 0 0 $X=18100 $Y=71950
X499 14 M2_M1_CDNS_7656752519023 $T=18260 81230 0 0 $X=18130 $Y=81150
X500 89 M2_M1_CDNS_7656752519023 $T=18960 81490 0 0 $X=18830 $Y=81410
X501 69 M2_M1_CDNS_7656752519023 $T=20130 89330 0 0 $X=20000 $Y=89250
X502 35 M2_M1_CDNS_7656752519023 $T=20130 103160 0 0 $X=20000 $Y=103080
X503 67 M2_M1_CDNS_7656752519023 $T=20370 44250 0 0 $X=20240 $Y=44170
X504 55 M2_M1_CDNS_7656752519023 $T=20550 72330 0 0 $X=20420 $Y=72250
X505 89 M2_M1_CDNS_7656752519023 $T=22920 81490 0 0 $X=22790 $Y=81410
X506 89 M2_M1_CDNS_7656752519023 $T=22920 82090 0 0 $X=22790 $Y=82010
X507 116 M2_M1_CDNS_7656752519023 $T=24280 44200 0 0 $X=24150 $Y=44120
X508 119 M2_M1_CDNS_7656752519023 $T=24390 101500 0 0 $X=24260 $Y=101420
X509 23 M2_M1_CDNS_7656752519023 $T=25170 80000 0 0 $X=25040 $Y=79920
X510 27 M2_M1_CDNS_7656752519023 $T=25170 97280 0 0 $X=25040 $Y=97200
X511 123 M2_M1_CDNS_7656752519023 $T=25890 64850 0 0 $X=25760 $Y=64770
X512 122 M2_M1_CDNS_7656752519023 $T=25910 72030 0 0 $X=25780 $Y=71950
X513 28 M2_M1_CDNS_7656752519023 $T=25910 97510 0 0 $X=25780 $Y=97430
X514 124 M2_M1_CDNS_7656752519023 $T=28230 72030 0 0 $X=28100 $Y=71950
X515 90 M2_M1_CDNS_7656752519023 $T=28230 79400 0 0 $X=28100 $Y=79320
X516 92 M2_M1_CDNS_7656752519023 $T=28230 89330 0 0 $X=28100 $Y=89250
X517 125 M2_M1_CDNS_7656752519023 $T=29570 73370 0 0 $X=29440 $Y=73290
X518 126 M2_M1_CDNS_7656752519023 $T=29570 81860 0 0 $X=29440 $Y=81780
X519 57 M2_M1_CDNS_7656752519023 $T=29570 90030 0 0 $X=29440 $Y=89950
X520 19 M2_M1_CDNS_7656752519023 $T=30510 99330 0 0 $X=30380 $Y=99250
X521 45 M2_M1_CDNS_7656752519023 $T=31430 100680 0 0 $X=31300 $Y=100600
X522 124 M2_M1_CDNS_7656752519023 $T=31890 72030 0 0 $X=31760 $Y=71950
X523 70 M2_M1_CDNS_7656752519023 $T=31890 98160 0 0 $X=31760 $Y=98080
X524 82 M2_M1_CDNS_7656752519023 $T=32630 73020 0 0 $X=32500 $Y=72940
X525 106 M2_M1_CDNS_7656752519023 $T=32630 97180 0 0 $X=32500 $Y=97100
X526 117 M2_M1_CDNS_7656752519023 $T=34080 44250 0 0 $X=33950 $Y=44170
X527 32 M2_M1_CDNS_7656752519023 $T=34650 101460 0 0 $X=34520 $Y=101380
X528 125 M2_M1_CDNS_7656752519023 $T=35300 73370 0 0 $X=35170 $Y=73290
X529 54 M2_M1_CDNS_7656752519023 $T=35430 96890 0 0 $X=35300 $Y=96810
X530 53 M2_M1_CDNS_7656752519023 $T=35830 97110 0 0 $X=35700 $Y=97030
X531 75 M2_M1_CDNS_7656752519023 $T=36510 80900 0 0 $X=36380 $Y=80820
X532 126 M2_M1_CDNS_7656752519023 $T=37250 81860 0 0 $X=37120 $Y=81780
X533 127 M2_M1_CDNS_7656752519023 $T=39570 72030 0 0 $X=39440 $Y=71950
X534 96 M2_M1_CDNS_7656752519023 $T=39570 81310 0 0 $X=39440 $Y=81230
X535 100 M2_M1_CDNS_7656752519023 $T=40910 72330 0 0 $X=40780 $Y=72250
X536 91 M2_M1_CDNS_7656752519023 $T=41210 98510 0 0 $X=41080 $Y=98430
X537 127 M2_M1_CDNS_7656752519023 $T=43230 72030 0 0 $X=43100 $Y=71950
X538 93 M2_M1_CDNS_7656752519023 $T=43230 89330 0 0 $X=43100 $Y=89250
X539 8 M2_M1_CDNS_7656752519023 $T=43920 101480 0 0 $X=43790 $Y=101400
X540 86 M2_M1_CDNS_7656752519023 $T=43970 71590 0 0 $X=43840 $Y=71510
X541 121 M2_M1_CDNS_7656752519023 $T=43970 80300 0 0 $X=43840 $Y=80220
X542 98 M2_M1_CDNS_7656752519023 $T=43970 98920 0 0 $X=43840 $Y=98840
X543 16 M2_M1_CDNS_7656752519023 $T=44250 100050 0 0 $X=44120 $Y=99970
X544 61 M2_M1_CDNS_7656752519023 $T=46480 100080 0 0 $X=46350 $Y=100000
X545 56 M2_M1_CDNS_7656752519023 $T=47850 80600 0 0 $X=47720 $Y=80520
X546 34 M2_M1_CDNS_7656752519023 $T=47850 88570 0 0 $X=47720 $Y=88490
X547 128 M2_M1_CDNS_7656752519023 $T=47980 64630 0 0 $X=47850 $Y=64550
X548 95 M2_M1_CDNS_7656752519023 $T=48590 90200 0 0 $X=48460 $Y=90120
X549 102 M2_M1_CDNS_7656752519023 $T=48600 99300 0 0 $X=48470 $Y=99220
X550 27 M2_M1_CDNS_7656752519023 $T=49320 99840 0 0 $X=49190 $Y=99760
X551 110 M2_M1_CDNS_7656752519023 $T=51270 96980 0 0 $X=51140 $Y=96900
X552 98 M2_M1_CDNS_7656752519023 $T=51700 98920 0 0 $X=51570 $Y=98840
X553 104 M2_M1_CDNS_7656752519023 $T=51940 82090 0 0 $X=51810 $Y=82010
X554 111 M2_M1_CDNS_7656752519023 $T=53770 97030 0 0 $X=53640 $Y=96950
X555 129 M2_M1_CDNS_7656752519023 $T=54180 98860 0 0 $X=54050 $Y=98780
X556 129 M2_M1_CDNS_7656752519023 $T=54180 100120 0 0 $X=54050 $Y=100040
X557 130 M2_M1_CDNS_7656752519023 $T=55000 97030 0 0 $X=54870 $Y=96950
X558 112 M2_M1_CDNS_7656752519023 $T=55250 73700 0 0 $X=55120 $Y=73620
X559 103 M2_M1_CDNS_7656752519023 $T=55290 71610 0 0 $X=55160 $Y=71530
X560 70 M2_M1_CDNS_7656752519023 $T=57720 100570 0 0 $X=57590 $Y=100490
X561 113 M2_M1_CDNS_7656752519023 $T=58070 101400 0 0 $X=57940 $Y=101320
X562 109 M2_M1_CDNS_7656752519023 $T=59200 80850 0 0 $X=59070 $Y=80770
X563 131 M2_M1_CDNS_7656752519023 $T=59410 91250 0 0 $X=59280 $Y=91170
X564 130 M2_M1_CDNS_7656752519023 $T=61910 97030 0 0 $X=61780 $Y=96950
X565 132 M2_M1_CDNS_7656752519025 $T=-260 63930 0 0 $X=-390 $Y=63800
X566 133 M2_M1_CDNS_7656752519025 $T=3160 97850 0 0 $X=3030 $Y=97720
X567 66 M2_M1_CDNS_7656752519025 $T=4450 38430 0 0 $X=4320 $Y=38300
X568 132 M2_M1_CDNS_7656752519025 $T=6890 63930 0 0 $X=6760 $Y=63800
X569 77 M2_M1_CDNS_7656752519025 $T=12420 38430 0 0 $X=12290 $Y=38300
X570 134 M2_M1_CDNS_7656752519025 $T=12890 59630 0 0 $X=12760 $Y=59500
X571 134 M2_M1_CDNS_7656752519025 $T=12890 64360 0 0 $X=12760 $Y=64230
X572 135 M2_M1_CDNS_7656752519025 $T=18230 63930 0 0 $X=18100 $Y=63800
X573 76 M2_M1_CDNS_7656752519025 $T=18990 38020 0 0 $X=18860 $Y=37890
X574 136 M2_M1_CDNS_7656752519025 $T=20570 64300 0 0 $X=20440 $Y=64170
X575 40 M2_M1_CDNS_7656752519025 $T=21290 80000 0 0 $X=21160 $Y=79870
X576 137 M2_M1_CDNS_7656752519025 $T=27340 60270 0 0 $X=27210 $Y=60140
X577 138 M2_M1_CDNS_7656752519025 $T=28230 63930 0 0 $X=28100 $Y=63800
X578 1 M2_M1_CDNS_7656752519025 $T=30220 101440 0 0 $X=30090 $Y=101310
X579 115 M2_M1_CDNS_7656752519025 $T=30820 16520 0 0 $X=30690 $Y=16390
X580 138 M2_M1_CDNS_7656752519025 $T=30840 58920 0 0 $X=30710 $Y=58790
X581 139 M2_M1_CDNS_7656752519025 $T=31460 59570 0 0 $X=31330 $Y=59440
X582 140 M2_M1_CDNS_7656752519025 $T=31730 37970 0 0 $X=31600 $Y=37840
X583 141 M2_M1_CDNS_7656752519025 $T=31750 16520 0 0 $X=31620 $Y=16390
X584 142 M2_M1_CDNS_7656752519025 $T=37230 64630 0 0 $X=37100 $Y=64500
X585 65 M2_M1_CDNS_7656752519025 $T=40080 38370 0 0 $X=39950 $Y=38240
X586 143 M2_M1_CDNS_7656752519025 $T=40910 64630 0 0 $X=40780 $Y=64500
X587 116 M2_M1_CDNS_7656752519025 $T=43970 17230 0 0 $X=43840 $Y=17100
X588 144 M2_M1_CDNS_7656752519025 $T=45670 38370 0 0 $X=45540 $Y=38240
X589 38 M2_M1_CDNS_7656752519025 $T=50120 100740 0 0 $X=49990 $Y=100610
X590 145 M2_M1_CDNS_7656752519025 $T=53980 60150 0 0 $X=53850 $Y=60020
X591 145 M2_M1_CDNS_7656752519025 $T=54640 63920 0 0 $X=54510 $Y=63790
X592 146 M2_M1_CDNS_7656752519025 $T=55250 65450 0 0 $X=55120 $Y=65320
X593 117 M2_M1_CDNS_7656752519025 $T=57490 16520 0 0 $X=57360 $Y=16390
X594 147 M2_M1_CDNS_7656752519025 $T=60810 32870 0 0 $X=60680 $Y=32740
X595 147 M2_M1_CDNS_7656752519025 $T=62710 101460 0 0 $X=62580 $Y=101330
X596 26 M3_M2_CDNS_7656752519026 $T=230 110810 0 0 $X=-20 $Y=110730
X597 3 M3_M2_CDNS_7656752519026 $T=20130 111380 0 0 $X=19880 $Y=111300
X598 39 M3_M2_CDNS_7656752519026 $T=21380 72640 0 0 $X=21130 $Y=72560
X599 28 M3_M2_CDNS_7656752519026 $T=25910 97510 0 0 $X=25660 $Y=97430
X600 115 M3_M2_CDNS_7656752519026 $T=30820 16520 0 0 $X=30570 $Y=16440
X601 138 M3_M2_CDNS_7656752519026 $T=30840 58920 0 0 $X=30590 $Y=58840
X602 141 M3_M2_CDNS_7656752519026 $T=31750 16520 0 0 $X=31500 $Y=16440
X603 65 M3_M2_CDNS_7656752519026 $T=59210 74060 0 0 $X=58960 $Y=73980
X604 144 M3_M2_CDNS_7656752519026 $T=59230 82660 0 0 $X=58980 $Y=82580
X605 140 M3_M2_CDNS_7656752519026 $T=59260 64440 0 0 $X=59010 $Y=64360
X606 47 M3_M2_CDNS_7656752519027 $T=550 64640 0 0 $X=470 $Y=64390
X607 87 M3_M2_CDNS_7656752519027 $T=2490 44290 0 0 $X=2410 $Y=44040
X608 12 M3_M2_CDNS_7656752519027 $T=2770 110920 0 0 $X=2690 $Y=110670
X609 74 M3_M2_CDNS_7656752519027 $T=7560 120840 0 0 $X=7480 $Y=120590
X610 47 M3_M2_CDNS_7656752519027 $T=11890 64220 0 0 $X=11810 $Y=63970
X611 83 M3_M2_CDNS_7656752519027 $T=17660 71070 0 0 $X=17580 $Y=70820
X612 123 M3_M2_CDNS_7656752519027 $T=22820 59760 0 0 $X=22740 $Y=59510
X613 47 M3_M2_CDNS_7656752519027 $T=23230 64170 0 0 $X=23150 $Y=63920
X614 64 M3_M2_CDNS_7656752519027 $T=25170 89190 0 0 $X=25090 $Y=88940
X615 83 M3_M2_CDNS_7656752519027 $T=28770 71070 0 0 $X=28690 $Y=70820
X616 47 M3_M2_CDNS_7656752519027 $T=34450 64130 0 0 $X=34370 $Y=63880
X617 142 M3_M2_CDNS_7656752519027 $T=35130 59760 0 0 $X=35050 $Y=59510
X618 83 M3_M2_CDNS_7656752519027 $T=40330 79760 0 0 $X=40250 $Y=79510
X619 47 M3_M2_CDNS_7656752519027 $T=45910 64110 0 0 $X=45830 $Y=63860
X620 83 M3_M2_CDNS_7656752519027 $T=51490 79650 0 0 $X=51410 $Y=79400
X621 47 M3_M2_CDNS_7656752519027 $T=57250 64080 0 0 $X=57170 $Y=63830
X622 47 M3_M2_CDNS_7656752519027 $T=59270 49170 0 180 $X=59190 $Y=48920
X623 47 M2_M1_CDNS_7656752519028 $T=550 64640 0 0 $X=470 $Y=64390
X624 87 M2_M1_CDNS_7656752519028 $T=2490 44290 0 0 $X=2410 $Y=44040
X625 12 M2_M1_CDNS_7656752519028 $T=2770 110920 0 0 $X=2690 $Y=110670
X626 74 M2_M1_CDNS_7656752519028 $T=7560 120840 0 0 $X=7480 $Y=120590
X627 47 M2_M1_CDNS_7656752519028 $T=11890 64220 0 0 $X=11810 $Y=63970
X628 83 M2_M1_CDNS_7656752519028 $T=17660 71070 0 0 $X=17580 $Y=70820
X629 47 M2_M1_CDNS_7656752519028 $T=23230 64170 0 0 $X=23150 $Y=63920
X630 64 M2_M1_CDNS_7656752519028 $T=25170 89190 0 0 $X=25090 $Y=88940
X631 83 M2_M1_CDNS_7656752519028 $T=28770 71070 0 0 $X=28690 $Y=70820
X632 47 M2_M1_CDNS_7656752519028 $T=34450 64130 0 0 $X=34370 $Y=63880
X633 83 M2_M1_CDNS_7656752519028 $T=40330 79760 0 0 $X=40250 $Y=79510
X634 47 M2_M1_CDNS_7656752519028 $T=45910 64110 0 0 $X=45830 $Y=63860
X635 83 M2_M1_CDNS_7656752519028 $T=51490 79650 0 0 $X=51410 $Y=79400
X636 47 M2_M1_CDNS_7656752519028 $T=57250 64080 0 0 $X=57170 $Y=63830
X637 133 M3_M2_CDNS_7656752519029 $T=3790 97850 0 0 $X=3660 $Y=97720
X638 132 M3_M2_CDNS_7656752519029 $T=4810 63930 0 0 $X=4680 $Y=63800
X639 115 M3_M2_CDNS_7656752519029 $T=9400 28030 0 0 $X=9270 $Y=27900
X640 123 M3_M2_CDNS_7656752519029 $T=22020 62580 0 0 $X=21890 $Y=62450
X641 76 M3_M2_CDNS_7656752519029 $T=25460 38020 0 0 $X=25330 $Y=37890
X642 76 M3_M2_CDNS_7656752519029 $T=28100 46420 0 0 $X=27970 $Y=46290
X643 78 M3_M2_CDNS_7656752519029 $T=31110 38400 0 0 $X=30980 $Y=38270
X644 139 M3_M2_CDNS_7656752519029 $T=31460 59570 0 0 $X=31330 $Y=59440
X645 142 M3_M2_CDNS_7656752519029 $T=37240 63760 0 0 $X=37110 $Y=63630
X646 117 M3_M2_CDNS_7656752519029 $T=57490 16820 0 0 $X=57360 $Y=16690
X647 14 M4_M3_CDNS_7656752519030 $T=6790 89980 0 0 $X=6420 $Y=89850
X648 25 M4_M3_CDNS_7656752519030 $T=9950 90030 0 0 $X=9580 $Y=89900
X649 20 M4_M3_CDNS_7656752519030 $T=37310 88780 0 0 $X=36940 $Y=88650
X650 27 M4_M3_CDNS_7656752519030 $T=49320 97160 0 0 $X=48950 $Y=97030
X651 71 M3_M2_CDNS_7656752519031 $T=8420 80300 0 0 $X=8290 $Y=80170
X652 68 M3_M2_CDNS_7656752519031 $T=9710 73550 0 0 $X=9580 $Y=73420
X653 35 M3_M2_CDNS_7656752519031 $T=20130 103160 0 0 $X=20000 $Y=103030
X654 66 M3_M2_CDNS_7656752519031 $T=41470 44250 0 0 $X=41340 $Y=44120
X655 76 M3_M2_CDNS_7656752519031 $T=52320 44250 0 0 $X=52190 $Y=44120
X656 9 M3_M2_CDNS_7656752519031 $T=54300 101520 0 0 $X=54170 $Y=101390
X657 14 M3_M2_CDNS_7656752519034 $T=18260 81230 0 0 $X=17890 $Y=81150
X658 60 M3_M2_CDNS_7656752519034 $T=51300 101400 0 0 $X=50930 $Y=101320
X659 66 M3_M2_CDNS_7656752519035 $T=4820 42750 0 0 $X=4740 $Y=42500
X660 4 M3_M2_CDNS_7656752519035 $T=22580 119930 0 0 $X=22500 $Y=119680
X661 133 M4_M3_CDNS_7656752519036 $T=-1050 17310 0 0 $X=-1130 $Y=17060
X662 4 M4_M3_CDNS_7656752519036 $T=22580 119930 0 0 $X=22500 $Y=119680
X663 49 M4_M3_CDNS_7656752519036 $T=37450 101760 0 0 $X=37370 $Y=101510
X664 47 M4_M3_CDNS_7656752519036 $T=60710 26810 0 0 $X=60630 $Y=26560
X665 132 M2_M1_CDNS_7656752519037 $T=-260 57410 0 0 $X=-390 $Y=57280
X666 80 M2_M1_CDNS_7656752519037 $T=870 59200 0 0 $X=740 $Y=59070
X667 148 M2_M1_CDNS_7656752519037 $T=3920 58640 0 0 $X=3790 $Y=58510
X668 132 M2_M1_CDNS_7656752519037 $T=4740 58230 0 0 $X=4610 $Y=58100
X669 84 M2_M1_CDNS_7656752519037 $T=5230 120900 0 0 $X=5100 $Y=120770
X670 148 M2_M1_CDNS_7656752519037 $T=8460 64880 0 0 $X=8330 $Y=64750
X671 149 M2_M1_CDNS_7656752519037 $T=12450 59070 0 0 $X=12320 $Y=58940
X672 149 M2_M1_CDNS_7656752519037 $T=12450 64880 0 0 $X=12320 $Y=64750
X673 133 M2_M1_CDNS_7656752519037 $T=13290 17310 0 0 $X=13160 $Y=17180
X674 39 M2_M1_CDNS_7656752519037 $T=13680 120910 0 0 $X=13550 $Y=120780
X675 136 M2_M1_CDNS_7656752519037 $T=17350 59970 0 0 $X=17220 $Y=59840
X676 135 M2_M1_CDNS_7656752519037 $T=18880 60150 0 0 $X=18750 $Y=60020
X677 123 M2_M1_CDNS_7656752519037 $T=22820 59760 0 0 $X=22690 $Y=59630
X678 137 M2_M1_CDNS_7656752519037 $T=30540 64940 0 0 $X=30410 $Y=64810
X679 78 M2_M1_CDNS_7656752519037 $T=31110 37850 0 0 $X=30980 $Y=37720
X680 139 M2_M1_CDNS_7656752519037 $T=31500 64270 0 0 $X=31370 $Y=64140
X681 142 M2_M1_CDNS_7656752519037 $T=35130 59760 0 0 $X=35000 $Y=59630
X682 67 M2_M1_CDNS_7656752519037 $T=37300 17230 0 0 $X=37170 $Y=17100
X683 150 M2_M1_CDNS_7656752519037 $T=39570 59570 0 0 $X=39440 $Y=59440
X684 150 M2_M1_CDNS_7656752519037 $T=39570 64630 0 0 $X=39440 $Y=64500
X685 66 M2_M1_CDNS_7656752519037 $T=41470 44250 0 0 $X=41340 $Y=44120
X686 97 M2_M1_CDNS_7656752519037 $T=43940 59990 0 0 $X=43810 $Y=59860
X687 143 M2_M1_CDNS_7656752519037 $T=45450 59630 0 0 $X=45320 $Y=59500
X688 77 M2_M1_CDNS_7656752519037 $T=46810 44250 0 0 $X=46680 $Y=44120
X689 101 M2_M1_CDNS_7656752519037 $T=49530 60010 0 0 $X=49400 $Y=59880
X690 76 M2_M1_CDNS_7656752519037 $T=52320 44250 0 0 $X=52190 $Y=44120
X691 78 M2_M1_CDNS_7656752519037 $T=54600 51480 0 0 $X=54470 $Y=51350
X692 131 M2_M1_CDNS_7656752519037 $T=58030 38310 0 0 $X=57900 $Y=38180
X693 128 M2_M1_CDNS_7656752519037 $T=58030 60140 0 0 $X=57900 $Y=60010
X694 146 M2_M1_CDNS_7656752519037 $T=60780 52610 0 0 $X=60650 $Y=52480
X695 151 M2_M1_CDNS_7656752519037 $T=61140 51440 0 0 $X=61010 $Y=51310
X696 151 M2_M1_CDNS_7656752519037 $T=61140 65420 0 0 $X=61010 $Y=65290
X697 115 M3_M2_CDNS_7656752519038 $T=-810 43780 0 0 $X=-940 $Y=43650
X698 141 M3_M2_CDNS_7656752519038 $T=-380 43220 0 0 $X=-510 $Y=43090
X699 115 M3_M2_CDNS_7656752519038 $T=10160 46120 0 0 $X=10030 $Y=45990
X700 77 M3_M2_CDNS_7656752519038 $T=12420 42300 0 0 $X=12290 $Y=42170
X701 67 M3_M2_CDNS_7656752519038 $T=22920 44250 0 0 $X=22790 $Y=44120
X702 66 M3_M2_CDNS_7656752519038 $T=27530 43890 0 0 $X=27400 $Y=43760
X703 138 M3_M2_CDNS_7656752519038 $T=31050 62810 0 0 $X=30920 $Y=62680
X704 78 M3_M2_CDNS_7656752519038 $T=31060 42750 0 0 $X=30930 $Y=42620
X705 139 M3_M2_CDNS_7656752519038 $T=31500 63160 0 0 $X=31370 $Y=63030
X706 140 M3_M2_CDNS_7656752519038 $T=31510 37970 0 0 $X=31380 $Y=37840
X707 141 M3_M2_CDNS_7656752519038 $T=31750 25000 0 0 $X=31620 $Y=24870
X708 65 M3_M2_CDNS_7656752519038 $T=40300 37320 0 0 $X=40170 $Y=37190
X709 144 M3_M2_CDNS_7656752519038 $T=45890 36750 0 0 $X=45760 $Y=36620
X710 77 M3_M2_CDNS_7656752519038 $T=46510 42300 0 0 $X=46380 $Y=42170
X711 117 M3_M2_CDNS_7656752519038 $T=50040 42300 0 0 $X=49910 $Y=42170
X712 117 M3_M2_CDNS_7656752519038 $T=50040 44310 0 0 $X=49910 $Y=44180
X713 78 M3_M2_CDNS_7656752519038 $T=54600 47040 0 0 $X=54470 $Y=46910
X714 78 M3_M2_CDNS_7656752519038 $T=55330 42750 0 0 $X=55200 $Y=42620
X715 65 M2_M1_CDNS_7656752519042 $T=59210 74060 0 0 $X=58960 $Y=73980
X716 144 M2_M1_CDNS_7656752519042 $T=59230 82660 0 0 $X=58980 $Y=82580
X717 77 M3_M2_CDNS_7656752519043 $T=13070 42750 0 0 $X=12820 $Y=42620
X718 76 M3_M2_CDNS_7656752519043 $T=18650 42750 0 0 $X=18400 $Y=42620
X719 77 M4_M3_CDNS_7656752519044 $T=13070 42750 0 0 $X=12820 $Y=42670
X720 116 M4_M3_CDNS_7656752519044 $T=61670 21020 0 0 $X=61420 $Y=20940
X721 117 M4_M3_CDNS_7656752519044 $T=62140 17310 0 0 $X=61890 $Y=17230
X722 66 M5_M4_CDNS_7656752519045 $T=4820 42750 0 0 $X=4740 $Y=42500
X723 65 M5_M4_CDNS_7656752519045 $T=40310 37330 0 0 $X=40230 $Y=37080
X724 67 M5_M4_CDNS_7656752519045 $T=60960 21490 0 0 $X=60880 $Y=21240
X725 65 M5_M4_CDNS_7656752519045 $T=61270 38260 0 0 $X=61190 $Y=38010
X726 67 M7_M6_CDNS_7656752519047 $T=22900 44330 0 0 $X=22770 $Y=44200
X727 116 M7_M6_CDNS_7656752519047 $T=27760 44330 0 0 $X=27630 $Y=44200
X728 116 M5_M4_CDNS_7656752519049 $T=61670 21020 0 0 $X=61420 $Y=20940
X729 117 M5_M4_CDNS_7656752519049 $T=62140 17310 0 0 $X=61890 $Y=17230
X730 116 M3_M2_CDNS_7656752519050 $T=61670 21020 0 0 $X=61420 $Y=20940
X731 117 M3_M2_CDNS_7656752519050 $T=62140 17310 0 0 $X=61890 $Y=17230
X732 67 M7_M6_CDNS_7656752519051 $T=60960 43450 0 0 $X=60830 $Y=43320
X733 116 M7_M6_CDNS_7656752519051 $T=61670 43980 0 0 $X=61540 $Y=43850
X734 117 M7_M6_CDNS_7656752519051 $T=62140 44330 0 0 $X=62010 $Y=44200
X735 116 M6_M5_CDNS_7656752519052 $T=61670 21020 0 0 $X=61420 $Y=20890
X736 117 M6_M5_CDNS_7656752519052 $T=62140 17310 0 0 $X=61890 $Y=17180
X737 67 M6_M5_CDNS_7656752519053 $T=60960 21490 0 0 $X=60880 $Y=21240
X738 133 M3_M2_CDNS_7656752519054 $T=-1050 17310 0 0 $X=-1180 $Y=17060
X739 67 M3_M2_CDNS_7656752519054 $T=60960 21490 0 0 $X=60830 $Y=21240
X740 133 M4_M3_CDNS_7656752519056 $T=3790 97120 0 0 $X=3660 $Y=96990
X741 116 M4_M3_CDNS_7656752519056 $T=22100 25350 0 0 $X=21970 $Y=25220
X742 117 M4_M3_CDNS_7656752519056 $T=57490 42300 0 0 $X=57360 $Y=42170
X743 116 M4_M3_CDNS_7656752519058 $T=18280 43890 0 0 $X=18150 $Y=43760
X744 78 M4_M3_CDNS_7656752519058 $T=54600 38400 0 0 $X=54470 $Y=38270
X745 117 M4_M3_CDNS_7656752519058 $T=57490 24370 0 0 $X=57360 $Y=24240
X746 115 M2_M1_CDNS_7656752519059 $T=7600 46120 0 0 $X=7470 $Y=45750
X747 141 M2_M1_CDNS_7656752519059 $T=15040 46000 0 0 $X=14910 $Y=45630
X748 65 M7_M6_CDNS_7656752519060 $T=40310 37330 0 0 $X=40230 $Y=37080
X749 65 M7_M6_CDNS_7656752519060 $T=61270 38260 0 0 $X=61190 $Y=38010
X750 65 M6_M5_CDNS_7656752519061 $T=40310 37330 0 0 $X=40230 $Y=37080
X751 65 M6_M5_CDNS_7656752519061 $T=61270 38260 0 0 $X=61190 $Y=38010
X752 118 47 79 10 48 83 241 240 600 809
+ 810 601 HAdder $T=-310 72840 0 0 $X=490 $Y=63880
X753 52 47 69 38 9 83 243 242 602 811
+ 812 603 HAdder $T=-310 98645 0 0 $X=490 $Y=89685
X754 80 47 133 79 119 83 245 244 604 813
+ 814 605 HAdder $T=-310 105415 0 0 $X=490 $Y=96455
X755 51 47 81 12 22 83 247 246 606 815
+ 816 607 HAdder $T=-310 112345 0 0 $X=490 $Y=103385
X756 120 47 152 84 32 83 249 248 608 817
+ 818 609 HAdder $T=12750 81440 1 180 $X=6160 $Y=72480
X757 55 47 153 74 51 83 251 250 610 819
+ 820 611 HAdder $T=11030 81440 0 0 $X=11830 $Y=72480
X758 121 47 86 85 154 83 253 252 612 821
+ 822 613 HAdder $T=11030 90040 0 0 $X=11830 $Y=81080
X759 34 47 56 11 46 83 255 254 614 823
+ 824 615 HAdder $T=24090 98645 1 180 $X=17500 $Y=89685
X760 128 47 101 155 100 83 257 256 616 825
+ 826 617 HAdder $T=45050 72840 0 0 $X=45850 $Y=63880
X761 146 47 145 156 103 83 259 258 618 827
+ 828 619 HAdder $T=58110 72840 1 180 $X=51520 $Y=63880
X762 112 47 156 107 104 83 261 260 620 829
+ 830 621 HAdder $T=58110 81440 1 180 $X=51520 $Y=72480
X763 140 47 151 157 112 83 263 262 622 831
+ 832 623 HAdder $T=56390 72840 0 0 $X=57190 $Y=63880
X764 65 47 157 158 109 83 265 264 624 833
+ 834 625 HAdder $T=56390 81440 0 0 $X=57190 $Y=72480
X765 144 47 158 159 114 83 267 266 626 835
+ 836 627 HAdder $T=56390 90040 0 0 $X=57190 $Y=81080
X766 131 47 159 160 113 83 269 268 628 837
+ 838 629 HAdder $T=56390 98640 0 0 $X=57190 $Y=89680
X767 87 132 80 148 47 83 115 149 134 141
+ 135 136 67 123 116 138 137 139 142 117
+ 66 150 97 77 143 101 76 128 145 78
+ 146 151 273 281 285 283 280 309 313 311
+ 308 270 287 291 296 279 315 319 324 272
+ 274 277 278 302 304 305 306 307 WallaceFinalAdder $T=0 42440 0 0 $X=0 $Y=42440
X768 47 71 45 82 50 161 83 334 333 332 FAdder $T=-600 81940 1 0 $X=490 $Y=72480
X769 47 42 41 161 13 36 83 337 336 335 FAdder $T=-600 90540 1 0 $X=490 $Y=81080
X770 47 162 21 163 26 81 83 340 339 338 FAdder $T=-600 109815 0 0 $X=490 $Y=110675
X771 47 132 152 148 68 118 83 343 342 341 FAdder $T=13040 73340 0 180 $X=6160 $Y=63880
X772 47 75 15 58 25 164 83 346 345 344 FAdder $T=13040 90540 0 180 $X=6160 $Y=81080
X773 47 73 43 164 30 16 83 349 348 347 FAdder $T=13040 99145 0 180 $X=6160 $Y=89685
X774 47 14 17 165 54 8 83 352 351 350 FAdder $T=13040 102525 1 180 $X=6160 $Y=103385
X775 47 166 1 167 18 165 83 355 354 353 FAdder $T=13040 109815 1 180 $X=6160 $Y=110675
X776 47 134 153 149 44 120 83 358 357 356 FAdder $T=10740 73340 1 0 $X=11830 $Y=63880
X777 47 20 5 154 49 24 83 361 360 359 FAdder $T=10740 99145 1 0 $X=11830 $Y=89685
X778 47 2 33 168 53 7 83 364 363 362 FAdder $T=10740 102525 0 0 $X=11830 $Y=103385
X779 47 169 19 170 29 168 83 367 366 365 FAdder $T=10740 109815 0 0 $X=11830 $Y=110675
X780 47 135 171 136 39 55 83 370 369 368 FAdder $T=24380 73340 0 180 $X=17500 $Y=63880
X781 47 122 172 171 40 14 83 373 372 371 FAdder $T=24380 81940 0 180 $X=17500 $Y=72480
X782 47 89 69 172 2 61 83 376 375 374 FAdder $T=24380 90540 0 180 $X=17500 $Y=81080
X783 47 64 35 173 59 6 83 379 378 377 FAdder $T=24380 102525 1 180 $X=17500 $Y=103385
X784 47 174 3 175 88 173 83 382 381 380 FAdder $T=24380 109815 1 180 $X=17500 $Y=110675
X785 47 138 176 123 4 122 83 385 384 383 FAdder $T=22080 73340 1 0 $X=23170 $Y=63880
X786 47 124 177 176 23 89 83 388 387 386 FAdder $T=22080 81940 1 0 $X=23170 $Y=72480
X787 47 90 178 177 64 52 83 391 390 389 FAdder $T=22080 90540 1 0 $X=23170 $Y=81080
X788 47 92 31 178 27 28 83 394 393 392 FAdder $T=22080 99145 1 0 $X=23170 $Y=89685
X789 47 139 179 137 82 124 83 397 396 395 FAdder $T=35720 73340 0 180 $X=28840 $Y=63880
X790 47 125 180 179 71 90 83 400 399 398 FAdder $T=35720 81940 0 180 $X=28840 $Y=72480
X791 47 126 181 180 42 92 83 403 402 401 FAdder $T=35720 90540 0 180 $X=28840 $Y=81080
X792 47 57 91 181 106 70 83 406 405 404 FAdder $T=35720 99145 0 180 $X=28840 $Y=89685
X793 47 150 182 142 58 125 83 409 408 407 FAdder $T=33420 73340 1 0 $X=34510 $Y=63880
X794 47 127 183 182 75 126 83 412 411 410 FAdder $T=33420 81940 1 0 $X=34510 $Y=72480
X795 47 96 184 183 73 57 83 415 414 413 FAdder $T=33420 90540 1 0 $X=34510 $Y=81080
X796 47 93 72 184 60 63 83 418 417 416 FAdder $T=33420 99145 1 0 $X=34510 $Y=89685
X797 47 143 185 97 86 127 83 421 420 419 FAdder $T=47060 73340 0 180 $X=40180 $Y=63880
X798 47 100 186 185 121 96 83 424 423 422 FAdder $T=47060 81940 0 180 $X=40180 $Y=72480
X799 47 94 187 186 20 93 83 427 426 425 FAdder $T=47060 90540 0 180 $X=40180 $Y=81080
X800 47 95 108 187 98 37 83 430 429 428 FAdder $T=47060 99145 0 180 $X=40180 $Y=89685
X801 47 103 188 155 56 94 83 433 432 431 FAdder $T=44760 81940 1 0 $X=45850 $Y=72480
X802 47 104 189 188 34 95 83 436 435 434 FAdder $T=44760 90540 1 0 $X=45850 $Y=81080
X803 47 105 110 189 99 102 83 439 438 437 FAdder $T=44760 99145 1 0 $X=45850 $Y=89685
X804 47 109 190 107 62 105 83 442 441 440 FAdder $T=58400 90540 0 180 $X=51520 $Y=81080
X805 47 114 111 190 129 130 83 445 444 443 FAdder $T=58400 99140 0 180 $X=51520 $Y=89680
X806 191 192 193 194 195 196 197 198 199 83
+ 37 102 130 160 147 47 28 70 63 200
+ 110 111 113 9 31 91 72 108 201 129
+ 38 27 106 60 98 99 202 61 36 16
+ 24 46 62 203 8 7 6 41 43 5
+ 11 22 17 33 35 204 13 30 49 32
+ 12 54 53 59 205 85 21 1 19 3
+ 45 15 206 48 18 29 88 50 25 119
+ 10 26 WallaceMultiplier $T=67110 70770 1 180 $X=23170 $Y=101330
X807 47 163 83 68 510 Diver $T=4340 118060 1 90 $X=490 $Y=118790
X808 47 162 83 84 511 Diver $T=7320 118060 1 90 $X=3470 $Y=118790
X809 47 166 83 74 512 Diver $T=5120 118010 0 90 $X=6160 $Y=118740
X810 47 167 83 44 513 Diver $T=8100 118050 0 90 $X=9140 $Y=118780
X811 47 170 83 39 514 Diver $T=15680 118090 1 90 $X=11830 $Y=118820
X812 47 169 83 40 515 Diver $T=18660 118080 1 90 $X=14810 $Y=118810
X813 47 174 83 23 516 Diver $T=16460 118040 0 90 $X=17500 $Y=118770
X814 47 175 83 4 517 Diver $T=19440 118020 0 90 $X=20480 $Y=118750
X815 207 66 47 83 208 209 210 211 212 133
+ 77 213 214 215 216 87 76 217 218 219
+ 220 78 115 141 140 221 222 223 224 225
+ 226 227 228 67 65 116 144 229 230 231
+ 232 233 234 235 117 131 236 237 238 147
+ 239 518 523 535 540 539 537 536 534 533
+ 572 571 578 577 574 573 570 542 548 547
+ 554 553 532 531 580 579 586 585 592 591
+ 521 525 524 528 527 530 529 562 561 564
+ 563 566 565 568 567 569 541 522 742 MAC $T=0 20 0 0 $X=0 $Y=20
M0 510 163 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=1270 $Y=119400 $dt=0
M1 68 510 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=1270 $Y=120330 $dt=0
M2 82 332 45 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=73900 $dt=0
M3 71 332 161 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=75240 $dt=0
M4 332 161 71 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=75650 $dt=0
M5 334 45 333 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=76580 $dt=0
M6 45 333 334 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=76990 $dt=0
M7 332 50 45 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=77400 $dt=0
M8 50 45 332 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=77810 $dt=0
M9 161 335 41 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=82500 $dt=0
M10 42 335 36 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=83840 $dt=0
M11 335 36 42 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=84250 $dt=0
M12 337 41 336 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=85180 $dt=0
M13 41 336 337 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=85590 $dt=0
M14 335 13 41 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=86000 $dt=0
M15 13 41 335 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=86410 $dt=0
M16 338 21 26 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=113855 $dt=0
M17 21 26 338 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=114265 $dt=0
M18 340 339 21 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=114675 $dt=0
M19 339 21 340 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=115085 $dt=0
M20 162 81 338 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=116015 $dt=0
M21 81 338 162 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=116425 $dt=0
M22 21 338 163 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=117765 $dt=0
M23 511 162 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=4250 $Y=119400 $dt=0
M24 84 511 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=4250 $Y=120330 $dt=0
M25 512 166 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=7950 $Y=119350 $dt=0
M26 74 512 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=7950 $Y=120280 $dt=0
M27 148 341 152 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=65300 $dt=0
M28 132 341 118 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=66640 $dt=0
M29 341 118 132 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=67050 $dt=0
M30 343 152 342 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=67980 $dt=0
M31 152 342 343 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=68390 $dt=0
M32 341 68 152 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=68800 $dt=0
M33 68 152 341 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=69210 $dt=0
M34 58 344 15 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=82500 $dt=0
M35 75 344 164 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=83840 $dt=0
M36 344 164 75 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=84250 $dt=0
M37 346 15 345 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=85180 $dt=0
M38 15 345 346 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=85590 $dt=0
M39 344 25 15 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=86000 $dt=0
M40 25 15 344 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=86410 $dt=0
M41 164 347 43 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=91105 $dt=0
M42 73 347 16 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=92445 $dt=0
M43 347 16 73 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=92855 $dt=0
M44 349 43 348 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=93785 $dt=0
M45 43 348 349 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=94195 $dt=0
M46 347 30 43 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=94605 $dt=0
M47 30 43 347 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=95015 $dt=0
M48 350 17 54 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=106565 $dt=0
M49 17 54 350 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=106975 $dt=0
M50 352 351 17 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=107385 $dt=0
M51 351 17 352 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=107795 $dt=0
M52 14 8 350 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=108725 $dt=0
M53 8 350 14 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=109135 $dt=0
M54 17 350 165 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=110475 $dt=0
M55 353 1 18 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=113855 $dt=0
M56 1 18 353 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=114265 $dt=0
M57 355 354 1 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=114675 $dt=0
M58 354 1 355 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=115085 $dt=0
M59 166 165 353 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=116015 $dt=0
M60 165 353 166 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=116425 $dt=0
M61 1 353 167 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=117765 $dt=0
M62 513 167 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=10930 $Y=119390 $dt=0
M63 44 513 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=10930 $Y=120320 $dt=0
M64 514 170 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=12610 $Y=119430 $dt=0
M65 39 514 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=12610 $Y=120360 $dt=0
M66 149 356 153 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=65300 $dt=0
M67 134 356 120 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=66640 $dt=0
M68 356 120 134 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=67050 $dt=0
M69 358 153 357 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=67980 $dt=0
M70 153 357 358 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=68390 $dt=0
M71 356 44 153 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=68800 $dt=0
M72 44 153 356 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=69210 $dt=0
M73 154 359 5 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=91105 $dt=0
M74 20 359 24 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=92445 $dt=0
M75 359 24 20 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=92855 $dt=0
M76 361 5 360 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=93785 $dt=0
M77 5 360 361 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=94195 $dt=0
M78 359 49 5 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=94605 $dt=0
M79 49 5 359 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=95015 $dt=0
M80 362 33 53 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=106565 $dt=0
M81 33 53 362 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=106975 $dt=0
M82 364 363 33 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=107385 $dt=0
M83 363 33 364 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=107795 $dt=0
M84 2 7 362 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=108725 $dt=0
M85 7 362 2 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=109135 $dt=0
M86 33 362 168 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=110475 $dt=0
M87 365 19 29 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=113855 $dt=0
M88 19 29 365 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=114265 $dt=0
M89 367 366 19 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=114675 $dt=0
M90 366 19 367 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=115085 $dt=0
M91 169 168 365 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=116015 $dt=0
M92 168 365 169 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=116425 $dt=0
M93 19 365 170 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=117765 $dt=0
M94 515 169 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=15590 $Y=119420 $dt=0
M95 40 515 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=15590 $Y=120350 $dt=0
M96 516 174 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=19290 $Y=119380 $dt=0
M97 23 516 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=19290 $Y=120310 $dt=0
M98 136 368 171 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.10357 scb=0.000255666 scc=3.44804e-08 $X=22160 $Y=65300 $dt=0
M99 135 368 55 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=66640 $dt=0
M100 368 55 135 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=67050 $dt=0
M101 370 171 369 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=67980 $dt=0
M102 171 369 370 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=68390 $dt=0
M103 368 39 171 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=68800 $dt=0
M104 39 171 368 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=69210 $dt=0
M105 171 371 172 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=73900 $dt=0
M106 122 371 14 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=75240 $dt=0
M107 371 14 122 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=75650 $dt=0
M108 373 172 372 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=76580 $dt=0
M109 172 372 373 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=76990 $dt=0
M110 371 40 172 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=77400 $dt=0
M111 40 172 371 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=77810 $dt=0
M112 172 374 69 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=82500 $dt=0
M113 89 374 61 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=83840 $dt=0
M114 374 61 89 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=84250 $dt=0
M115 376 69 375 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=85180 $dt=0
M116 69 375 376 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=85590 $dt=0
M117 374 2 69 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=86000 $dt=0
M118 2 69 374 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=86410 $dt=0
M119 377 35 59 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=106565 $dt=0
M120 35 59 377 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=106975 $dt=0
M121 379 378 35 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=107385 $dt=0
M122 378 35 379 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=107795 $dt=0
M123 64 6 377 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=108725 $dt=0
M124 6 377 64 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=109135 $dt=0
M125 35 377 173 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=110475 $dt=0
M126 380 3 88 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=113855 $dt=0
M127 3 88 380 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=114265 $dt=0
M128 382 381 3 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=114675 $dt=0
M129 381 3 382 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=4.11282 scb=0.000306462 scc=1.0989e-07 $X=22160 $Y=115085 $dt=0
M130 174 173 380 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=116015 $dt=0
M131 173 380 174 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=116425 $dt=0
M132 3 380 175 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=117765 $dt=0
M133 517 175 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=22270 $Y=119360 $dt=0
M134 4 517 47 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8263 scb=0.00911451 scc=0.000207374 $X=22270 $Y=120290 $dt=0
M135 123 383 176 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=65300 $dt=0
M136 138 383 122 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=66640 $dt=0
M137 383 122 138 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=67050 $dt=0
M138 385 176 384 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=67980 $dt=0
M139 176 384 385 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=68390 $dt=0
M140 383 4 176 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=68800 $dt=0
M141 4 176 383 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=69210 $dt=0
M142 176 386 177 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=73900 $dt=0
M143 124 386 89 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=75240 $dt=0
M144 386 89 124 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=75650 $dt=0
M145 388 177 387 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=76580 $dt=0
M146 177 387 388 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=76990 $dt=0
M147 386 23 177 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=77400 $dt=0
M148 23 177 386 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=77810 $dt=0
M149 177 389 178 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=82500 $dt=0
M150 90 389 52 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=83840 $dt=0
M151 389 52 90 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=84250 $dt=0
M152 391 178 390 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=85180 $dt=0
M153 178 390 391 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=85590 $dt=0
M154 389 64 178 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=86000 $dt=0
M155 64 178 389 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=86410 $dt=0
M156 178 392 31 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=91105 $dt=0
M157 92 392 28 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=92445 $dt=0
M158 392 28 92 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=92855 $dt=0
M159 394 31 393 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=93785 $dt=0
M160 31 393 394 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=94195 $dt=0
M161 392 27 31 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=94605 $dt=0
M162 27 31 392 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=95015 $dt=0
M163 137 395 179 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.10624 scb=0.000256891 scc=3.49982e-08 $X=33500 $Y=65300 $dt=0
M164 139 395 124 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=66640 $dt=0
M165 395 124 139 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=67050 $dt=0
M166 397 179 396 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=67980 $dt=0
M167 179 396 397 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=68390 $dt=0
M168 395 82 179 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=68800 $dt=0
M169 82 179 395 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=69210 $dt=0
M170 179 398 180 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=73900 $dt=0
M171 125 398 90 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=75240 $dt=0
M172 398 90 125 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=75650 $dt=0
M173 400 180 399 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=76580 $dt=0
M174 180 399 400 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=76990 $dt=0
M175 398 71 180 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=77400 $dt=0
M176 71 180 398 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=77810 $dt=0
M177 180 401 181 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=82500 $dt=0
M178 126 401 92 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=83840 $dt=0
M179 401 92 126 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=84250 $dt=0
M180 403 181 402 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=85180 $dt=0
M181 181 402 403 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=85590 $dt=0
M182 401 42 181 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=86000 $dt=0
M183 42 181 401 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=86410 $dt=0
M184 181 404 91 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=91105 $dt=0
M185 57 404 70 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=92445 $dt=0
M186 404 70 57 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=92855 $dt=0
M187 406 91 405 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=93785 $dt=0
M188 91 405 406 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=94195 $dt=0
M189 404 106 91 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=94605 $dt=0
M190 106 91 404 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=95015 $dt=0
M191 142 407 182 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.71642 scb=0.000135303 scc=5.64513e-09 $X=35400 $Y=65300 $dt=0
M192 150 407 125 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=66640 $dt=0
M193 407 125 150 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=67050 $dt=0
M194 409 182 408 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=67980 $dt=0
M195 182 408 409 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=68390 $dt=0
M196 407 58 182 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=68800 $dt=0
M197 58 182 407 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=69210 $dt=0
M198 182 410 183 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=73900 $dt=0
M199 127 410 126 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=75240 $dt=0
M200 410 126 127 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=75650 $dt=0
M201 412 183 411 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=76580 $dt=0
M202 183 411 412 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=76990 $dt=0
M203 410 75 183 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=77400 $dt=0
M204 75 183 410 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=77810 $dt=0
M205 183 413 184 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=82500 $dt=0
M206 96 413 57 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=83840 $dt=0
M207 413 57 96 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=84250 $dt=0
M208 415 184 414 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=85180 $dt=0
M209 184 414 415 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=85590 $dt=0
M210 413 73 184 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=86000 $dt=0
M211 73 184 413 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=86410 $dt=0
M212 184 416 72 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=91105 $dt=0
M213 93 416 63 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=92445 $dt=0
M214 416 63 93 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=92855 $dt=0
M215 418 72 417 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=93785 $dt=0
M216 72 417 418 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=94195 $dt=0
M217 416 60 72 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=94605 $dt=0
M218 60 72 416 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=95015 $dt=0
M219 97 419 185 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=65300 $dt=0
M220 143 419 127 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=66640 $dt=0
M221 419 127 143 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=67050 $dt=0
M222 421 185 420 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=67980 $dt=0
M223 185 420 421 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=68390 $dt=0
M224 419 86 185 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=68800 $dt=0
M225 86 185 419 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=69210 $dt=0
M226 185 422 186 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=73900 $dt=0
M227 100 422 96 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=75240 $dt=0
M228 422 96 100 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=75650 $dt=0
M229 424 186 423 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=76580 $dt=0
M230 186 423 424 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=76990 $dt=0
M231 422 121 186 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=77400 $dt=0
M232 121 186 422 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=77810 $dt=0
M233 186 425 187 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=82500 $dt=0
M234 94 425 93 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=83840 $dt=0
M235 425 93 94 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=84250 $dt=0
M236 427 187 426 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=85180 $dt=0
M237 187 426 427 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=85590 $dt=0
M238 425 20 187 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=86000 $dt=0
M239 20 187 425 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=86410 $dt=0
M240 187 428 108 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=91105 $dt=0
M241 95 428 37 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=92445 $dt=0
M242 428 37 95 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=92855 $dt=0
M243 430 108 429 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=93785 $dt=0
M244 108 429 430 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=94195 $dt=0
M245 428 98 108 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=94605 $dt=0
M246 98 108 428 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=95015 $dt=0
M247 155 431 188 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=73900 $dt=0
M248 103 431 94 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=75240 $dt=0
M249 431 94 103 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=75650 $dt=0
M250 433 188 432 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=76580 $dt=0
M251 188 432 433 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=76990 $dt=0
M252 431 56 188 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=77400 $dt=0
M253 56 188 431 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=77810 $dt=0
M254 188 434 189 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=82500 $dt=0
M255 104 434 95 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=83840 $dt=0
M256 434 95 104 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=84250 $dt=0
M257 436 189 435 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=85180 $dt=0
M258 189 435 436 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=85590 $dt=0
M259 434 34 189 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=86000 $dt=0
M260 34 189 434 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=86410 $dt=0
M261 189 437 110 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=91105 $dt=0
M262 105 437 102 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=92445 $dt=0
M263 437 102 105 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=92855 $dt=0
M264 439 110 438 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=93785 $dt=0
M265 110 438 439 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=94195 $dt=0
M266 437 99 110 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=94605 $dt=0
M267 99 110 437 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=95015 $dt=0
M268 107 440 190 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=82500 $dt=0
M269 109 440 105 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=83840 $dt=0
M270 440 105 109 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=84250 $dt=0
M271 442 190 441 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=85180 $dt=0
M272 190 441 442 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=85590 $dt=0
M273 440 62 190 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=86000 $dt=0
M274 62 190 440 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=86410 $dt=0
M275 190 443 111 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=91100 $dt=0
M276 114 443 130 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=92440 $dt=0
M277 443 130 114 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=92850 $dt=0
M278 445 111 444 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=93780 $dt=0
M279 111 444 445 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=94190 $dt=0
M280 443 129 111 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=94600 $dt=0
M281 129 111 443 47 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=95010 $dt=0
M282 510 163 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=2280 $Y=119400 $dt=1
M283 68 510 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=2280 $Y=120330 $dt=1
M284 82 332 161 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=4830 $Y=73900 $dt=1
M285 161 335 36 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=4830 $Y=82500 $dt=1
M286 81 338 163 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=4830 $Y=117765 $dt=1
M287 810 241 79 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=65950 $dt=1
M288 83 240 810 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=5210 $Y=66160 $dt=1
M289 83 240 809 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=5210 $Y=67090 $dt=1
M290 809 241 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=5210 $Y=67500 $dt=1
M291 118 48 809 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=67910 $dt=1
M292 809 10 118 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=68320 $dt=1
M293 83 10 240 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5210 $Y=69250 $dt=1
M294 83 48 241 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=70180 $dt=1
M295 812 243 69 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=91755 $dt=1
M296 83 242 812 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=5210 $Y=91965 $dt=1
M297 83 242 811 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=5210 $Y=92895 $dt=1
M298 811 243 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=5210 $Y=93305 $dt=1
M299 52 9 811 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=93715 $dt=1
M300 811 38 52 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=94125 $dt=1
M301 83 38 242 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5210 $Y=95055 $dt=1
M302 83 9 243 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=95985 $dt=1
M303 814 245 133 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5210 $Y=98525 $dt=1
M304 83 244 814 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=5210 $Y=98735 $dt=1
M305 83 244 813 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=5210 $Y=99665 $dt=1
M306 813 245 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=5210 $Y=100075 $dt=1
M307 80 119 813 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=5210 $Y=100485 $dt=1
M308 813 79 80 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=5210 $Y=100895 $dt=1
M309 83 79 244 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=5210 $Y=101825 $dt=1
M310 83 119 245 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5210 $Y=102755 $dt=1
M311 816 247 81 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=105455 $dt=1
M312 83 246 816 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=5210 $Y=105665 $dt=1
M313 83 246 815 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=5210 $Y=106595 $dt=1
M314 815 247 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=5210 $Y=107005 $dt=1
M315 51 22 815 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=107415 $dt=1
M316 815 12 51 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=107825 $dt=1
M317 83 12 246 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5210 $Y=108755 $dt=1
M318 83 22 247 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=109685 $dt=1
M319 511 162 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=5260 $Y=119400 $dt=1
M320 84 511 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=5260 $Y=120330 $dt=1
M321 512 166 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=6940 $Y=119350 $dt=1
M322 74 512 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=6940 $Y=120280 $dt=1
M323 818 249 152 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=6990 $Y=74550 $dt=1
M324 83 248 818 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=6990 $Y=74760 $dt=1
M325 83 248 817 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=6990 $Y=75690 $dt=1
M326 817 249 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=6990 $Y=76100 $dt=1
M327 120 32 817 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6990 $Y=76510 $dt=1
M328 817 84 120 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6990 $Y=76920 $dt=1
M329 83 84 248 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=6990 $Y=77850 $dt=1
M330 83 32 249 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=6990 $Y=78780 $dt=1
M331 148 341 118 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=7370 $Y=65300 $dt=1
M332 58 344 164 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=7370 $Y=82500 $dt=1
M333 164 347 16 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=7370 $Y=91105 $dt=1
M334 8 350 165 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=7370 $Y=110475 $dt=1
M335 165 353 167 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=7370 $Y=117765 $dt=1
M336 513 167 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=9920 $Y=119390 $dt=1
M337 44 513 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=9920 $Y=120320 $dt=1
M338 514 170 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=13620 $Y=119430 $dt=1
M339 39 514 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=13620 $Y=120360 $dt=1
M340 149 356 120 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=16170 $Y=65300 $dt=1
M341 154 359 24 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=16170 $Y=91105 $dt=1
M342 7 362 168 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=16170 $Y=110475 $dt=1
M343 168 365 170 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=16170 $Y=117765 $dt=1
M344 820 251 153 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=74550 $dt=1
M345 83 250 820 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=16550 $Y=74760 $dt=1
M346 83 250 819 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=16550 $Y=75690 $dt=1
M347 819 251 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=16550 $Y=76100 $dt=1
M348 55 51 819 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=76510 $dt=1
M349 819 74 55 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=76920 $dt=1
M350 83 74 250 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=16550 $Y=77850 $dt=1
M351 83 51 251 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=78780 $dt=1
M352 822 253 86 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=83150 $dt=1
M353 83 252 822 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=16550 $Y=83360 $dt=1
M354 83 252 821 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=16550 $Y=84290 $dt=1
M355 821 253 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=16550 $Y=84700 $dt=1
M356 121 154 821 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=85110 $dt=1
M357 821 85 121 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=85520 $dt=1
M358 83 85 252 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=16550 $Y=86450 $dt=1
M359 83 154 253 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=87380 $dt=1
M360 515 169 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=16600 $Y=119420 $dt=1
M361 40 515 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=16600 $Y=120350 $dt=1
M362 516 174 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=18280 $Y=119380 $dt=1
M363 23 516 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=18280 $Y=120310 $dt=1
M364 824 255 56 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=18330 $Y=91755 $dt=1
M365 83 254 824 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=18330 $Y=91965 $dt=1
M366 83 254 823 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=18330 $Y=92895 $dt=1
M367 823 255 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=18330 $Y=93305 $dt=1
M368 34 46 823 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=18330 $Y=93715 $dt=1
M369 823 11 34 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=18330 $Y=94125 $dt=1
M370 83 11 254 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=18330 $Y=95055 $dt=1
M371 83 46 255 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=18330 $Y=95985 $dt=1
M372 136 368 55 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=18710 $Y=65300 $dt=1
M373 171 371 14 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=18710 $Y=73900 $dt=1
M374 172 374 61 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=18710 $Y=82500 $dt=1
M375 6 377 173 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=18710 $Y=110475 $dt=1
M376 173 380 175 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=18710 $Y=117765 $dt=1
M377 517 175 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=21260 $Y=119360 $dt=1
M378 4 517 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=21260 $Y=120290 $dt=1
M379 123 383 122 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=65300 $dt=1
M380 176 386 89 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=73900 $dt=1
M381 177 389 52 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=82500 $dt=1
M382 178 392 28 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=91105 $dt=1
M383 137 395 124 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=65300 $dt=1
M384 179 398 90 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=73900 $dt=1
M385 180 401 92 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=82500 $dt=1
M386 181 404 70 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=91105 $dt=1
M387 142 407 125 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=65300 $dt=1
M388 182 410 126 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=73900 $dt=1
M389 183 413 57 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=82500 $dt=1
M390 184 416 63 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=91105 $dt=1
M391 97 419 127 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=65300 $dt=1
M392 185 422 96 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=73900 $dt=1
M393 186 425 93 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=82500 $dt=1
M394 187 428 37 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=91105 $dt=1
M395 155 431 94 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=50190 $Y=73900 $dt=1
M396 188 434 95 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=50190 $Y=82500 $dt=1
M397 189 437 102 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=50190 $Y=91105 $dt=1
M398 826 257 101 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=50570 $Y=65950 $dt=1
M399 83 256 826 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.901 scb=0.0471116 scc=0.0116656 $X=50570 $Y=66160 $dt=1
M400 83 256 825 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.1268 scb=0.0349743 scc=0.0111863 $X=50570 $Y=67090 $dt=1
M401 825 257 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.5388 scb=0.0347327 scc=0.0111862 $X=50570 $Y=67500 $dt=1
M402 128 100 825 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=50570 $Y=67910 $dt=1
M403 825 155 128 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=50570 $Y=68320 $dt=1
M404 83 155 256 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.6513 scb=0.0354006 scc=0.011187 $X=50570 $Y=69250 $dt=1
M405 83 100 257 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=50570 $Y=70180 $dt=1
M406 828 259 145 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=52350 $Y=65950 $dt=1
M407 83 258 828 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.901 scb=0.0471116 scc=0.0116656 $X=52350 $Y=66160 $dt=1
M408 83 258 827 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.1268 scb=0.0349743 scc=0.0111863 $X=52350 $Y=67090 $dt=1
M409 827 259 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.5388 scb=0.0347327 scc=0.0111862 $X=52350 $Y=67500 $dt=1
M410 146 103 827 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=52350 $Y=67910 $dt=1
M411 827 156 146 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=52350 $Y=68320 $dt=1
M412 83 156 258 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.6513 scb=0.0354006 scc=0.011187 $X=52350 $Y=69250 $dt=1
M413 83 103 259 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=52350 $Y=70180 $dt=1
M414 830 261 156 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52350 $Y=74550 $dt=1
M415 83 260 830 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=52350 $Y=74760 $dt=1
M416 83 260 829 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=52350 $Y=75690 $dt=1
M417 829 261 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=52350 $Y=76100 $dt=1
M418 112 104 829 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52350 $Y=76510 $dt=1
M419 829 107 112 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52350 $Y=76920 $dt=1
M420 83 107 260 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=52350 $Y=77850 $dt=1
M421 83 104 261 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52350 $Y=78780 $dt=1
M422 107 440 105 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52730 $Y=82500 $dt=1
M423 190 443 130 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52730 $Y=91100 $dt=1
M424 832 263 151 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=65950 $dt=1
M425 83 262 832 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=66160 $dt=1
M426 83 262 831 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=67090 $dt=1
M427 831 263 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=67500 $dt=1
M428 140 112 831 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=67910 $dt=1
M429 831 157 140 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=68320 $dt=1
M430 83 157 262 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=69250 $dt=1
M431 83 112 263 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=70180 $dt=1
M432 834 265 157 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=74550 $dt=1
M433 83 264 834 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=74760 $dt=1
M434 83 264 833 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=75690 $dt=1
M435 833 265 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=76100 $dt=1
M436 65 109 833 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=76510 $dt=1
M437 833 158 65 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=76920 $dt=1
M438 83 158 264 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=77850 $dt=1
M439 83 109 265 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=78780 $dt=1
M440 836 267 158 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=83150 $dt=1
M441 83 266 836 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=83360 $dt=1
M442 83 266 835 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=84290 $dt=1
M443 835 267 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=84700 $dt=1
M444 144 114 835 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=85110 $dt=1
M445 835 159 144 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=85520 $dt=1
M446 83 159 266 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=86450 $dt=1
M447 83 114 267 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=87380 $dt=1
M448 838 269 159 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=91750 $dt=1
M449 83 268 838 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=91960 $dt=1
M450 83 268 837 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=92890 $dt=1
M451 837 269 83 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=93300 $dt=1
M452 131 113 837 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=93710 $dt=1
M453 837 160 131 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=94120 $dt=1
M454 83 160 268 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=95050 $dt=1
M455 83 113 269 83 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=95980 $dt=1
.ends WallaceProjectMAC
