* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : WallaceFinalAdder                            *
* Netlisted  : Thu Dec 11 09:02:36 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765461750680                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765461750680 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765461750680

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765461750681                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765461750681 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765461750681

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765461750682                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765461750682 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765461750682

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765461750683                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765461750683 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765461750683

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765461750684                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765461750684 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765461750684

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765461750685                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765461750685 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765461750685

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765461750686                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765461750686 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765461750686

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765461750687                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765461750687 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765461750687

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765461750688                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765461750688 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765461750688

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765461750689                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765461750689 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765461750689

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7654617506810                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7654617506810 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7654617506810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7654617506811                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7654617506811 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7654617506811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7654617506812                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7654617506812 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7654617506812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7654617506813                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7654617506813 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7654617506813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7654617506814                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7654617506814 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7654617506814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750680                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750680 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750680

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750681                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750681 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765461750681

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750682                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750682 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750682

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750683                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750683 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765461750683

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750684                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750684 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765461750684

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750685                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750685 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750685

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X0 1 M2_M1_CDNS_765461750683 $T=1510 -2070 0 0 $X=1430 $Y=-2200
X1 1 M2_M1_CDNS_765461750683 $T=3010 -2070 0 0 $X=2930 $Y=-2200
X2 2 M1_PO_CDNS_7654617506812 $T=1870 -1670 0 0 $X=1770 $Y=-1790
X3 1 M1_PO_CDNS_7654617506812 $T=2510 -2070 0 0 $X=2410 $Y=-2190
X4 6 M1_PO_CDNS_7654617506812 $T=4500 -2020 0 0 $X=4400 $Y=-2140
X5 5 M3_M2_CDNS_7654617506813 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X6 5 M2_M1_CDNS_7654617506814 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X7 4 5 6 nmos1v_CDNS_765461750680 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X8 3 5 6 4 pmos1v_CDNS_765461750681 $T=4560 -1510 0 0 $X=3880 $Y=-1710
X9 4 1 7 nmos1v_CDNS_765461750682 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X10 3 2 6 4 pmos1v_CDNS_765461750683 $T=1930 -1320 0 0 $X=1250 $Y=-1520
X11 3 6 1 4 pmos1v_CDNS_765461750684 $T=2430 -1320 1 180 $X=1980 $Y=-1520
X12 6 2 7 4 nmos1v_CDNS_765461750685 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7654617506815                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7654617506815 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7654617506815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7654617506816                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7654617506816 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7654617506816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750686                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750686 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765461750686

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750687                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750687 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750687

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X0 6 M2_M1_CDNS_765461750683 $T=690 3330 0 0 $X=610 $Y=3200
X1 1 M2_M1_CDNS_765461750683 $T=1190 1490 0 0 $X=1110 $Y=1360
X2 1 M2_M1_CDNS_765461750683 $T=2520 1490 0 0 $X=2440 $Y=1360
X3 6 M2_M1_CDNS_765461750683 $T=2550 3330 0 0 $X=2470 $Y=3200
X4 4 M5_M4_CDNS_765461750684 $T=1850 2810 0 90 $X=1600 $Y=2590
X5 4 M4_M3_CDNS_765461750686 $T=1850 2810 0 90 $X=1600 $Y=2590
X6 4 M3_M2_CDNS_765461750687 $T=1850 2810 0 90 $X=1600 $Y=2590
X7 4 M2_M1_CDNS_765461750688 $T=1850 2810 0 90 $X=1600 $Y=2590
X8 4 M6_M5_CDNS_765461750689 $T=1850 2810 0 90 $X=1600 $Y=2590
X9 7 M1_PO_CDNS_7654617506812 $T=2470 2570 0 0 $X=2370 $Y=2450
X10 1 M1_PO_CDNS_7654617506815 $T=320 1490 0 0 $X=220 $Y=1240
X11 5 M1_PO_CDNS_7654617506815 $T=1540 2050 0 0 $X=1440 $Y=1800
X12 5 M1_PO_CDNS_7654617506815 $T=3400 2050 0 0 $X=3300 $Y=1800
X13 1 M2_M1_CDNS_7654617506816 $T=320 1490 0 0 $X=240 $Y=1240
X14 5 M2_M1_CDNS_7654617506816 $T=1540 2050 0 0 $X=1460 $Y=1800
X15 5 M2_M1_CDNS_7654617506816 $T=3400 2050 0 0 $X=3320 $Y=1800
X16 2 2 1 6 3 pmos1v_CDNS_765461750686 $T=420 3660 0 0 $X=0 $Y=3460
X17 1 2 5 4 3 pmos1v_CDNS_765461750686 $T=1350 3660 0 0 $X=930 $Y=3460
X18 6 2 7 4 3 pmos1v_CDNS_765461750686 $T=2370 3660 1 180 $X=1860 $Y=3460
X19 2 2 5 7 3 pmos1v_CDNS_765461750686 $T=3300 3660 1 180 $X=2790 $Y=3460
X20 3 3 1 6 nmos1v_CDNS_765461750687 $T=420 800 0 0 $X=0 $Y=240
X21 4 3 5 6 nmos1v_CDNS_765461750687 $T=1440 800 1 180 $X=930 $Y=240
X22 4 3 7 1 nmos1v_CDNS_765461750687 $T=2280 800 0 0 $X=1860 $Y=240
X23 3 3 5 7 nmos1v_CDNS_765461750687 $T=3300 800 1 180 $X=2790 $Y=240
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7654617506818                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7654617506818 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7654617506818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7654617506819                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7654617506819 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7654617506819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7654617506820                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7654617506820 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7654617506820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750688                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750688 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765461750688

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750689                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750689 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750689

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506810                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506810 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506811                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506811 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506812                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506812 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506813                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506813 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7654617506813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506814                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506814 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506815                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506815 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506816                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506816 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506817                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506817 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506818                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506818 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=16
X0 1 M2_M1_CDNS_765461750683 $T=2220 -7390 0 90 $X=2090 $Y=-7470
X1 1 M2_M1_CDNS_765461750683 $T=2220 -4680 0 90 $X=2090 $Y=-4760
X2 7 M2_M1_CDNS_765461750683 $T=4200 -2840 0 90 $X=4070 $Y=-2920
X3 8 M2_M1_CDNS_765461750683 $T=4570 -3920 0 90 $X=4440 $Y=-4000
X4 8 M1_PO_CDNS_7654617506815 $T=2340 -4370 0 90 $X=2090 $Y=-4470
X5 8 M1_PO_CDNS_7654617506815 $T=2930 -6480 0 90 $X=2680 $Y=-6580
X6 8 M1_PO_CDNS_7654617506815 $T=2950 -5710 0 90 $X=2700 $Y=-5810
X7 4 M1_PO_CDNS_7654617506815 $T=3490 -4140 0 90 $X=3240 $Y=-4240
X8 4 M1_PO_CDNS_7654617506815 $T=3500 -3460 0 90 $X=3250 $Y=-3560
X9 8 M2_M1_CDNS_7654617506816 $T=2340 -4370 0 90 $X=2090 $Y=-4450
X10 8 M2_M1_CDNS_7654617506816 $T=2930 -6480 0 90 $X=2680 $Y=-6560
X11 8 M2_M1_CDNS_7654617506816 $T=2950 -5710 0 90 $X=2700 $Y=-5790
X12 4 M2_M1_CDNS_7654617506816 $T=3490 -4140 0 90 $X=3240 $Y=-4220
X13 4 M2_M1_CDNS_7654617506816 $T=3500 -3460 0 90 $X=3250 $Y=-3540
X14 9 M2_M1_CDNS_7654617506816 $T=5640 -5920 0 90 $X=5390 $Y=-6000
X15 9 M2_M1_CDNS_7654617506816 $T=5640 -5080 0 90 $X=5390 $Y=-5160
X16 9 M2_M1_CDNS_7654617506816 $T=5640 -4300 0 90 $X=5390 $Y=-4380
X17 6 6 4 8 2 pmos1v_CDNS_765461750686 $T=5520 -3500 0 270 $X=5320 $Y=-4010
X18 6 6 5 7 2 pmos1v_CDNS_765461750686 $T=5520 -2570 0 270 $X=5320 $Y=-3080
X19 2 2 4 8 nmos1v_CDNS_765461750687 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X20 2 2 5 7 nmos1v_CDNS_765461750687 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X21 10 M2_M1_CDNS_7654617506818 $T=1300 -5710 0 90 $X=1170 $Y=-5840
X22 10 M2_M1_CDNS_7654617506818 $T=1300 -4270 0 90 $X=1170 $Y=-4400
X23 4 M2_M1_CDNS_7654617506819 $T=3500 -4810 0 0 $X=3250 $Y=-4940
X24 4 M2_M1_CDNS_7654617506819 $T=3500 -1930 0 0 $X=3250 $Y=-2060
X25 7 M2_M1_CDNS_7654617506819 $T=4210 -6730 0 0 $X=3960 $Y=-6860
X26 7 M2_M1_CDNS_7654617506819 $T=4210 -5370 0 0 $X=3960 $Y=-5500
X27 8 M2_M1_CDNS_7654617506819 $T=4540 -5740 0 0 $X=4290 $Y=-5870
X28 5 M2_M1_CDNS_7654617506819 $T=4960 -4960 0 0 $X=4710 $Y=-5090
X29 5 M2_M1_CDNS_7654617506819 $T=4960 -2500 0 0 $X=4710 $Y=-2630
X30 4 M1_PO_CDNS_7654617506820 $T=3500 -4810 0 0 $X=3260 $Y=-4910
X31 7 M1_PO_CDNS_7654617506820 $T=4210 -6730 0 0 $X=3970 $Y=-6830
X32 7 M1_PO_CDNS_7654617506820 $T=4210 -5370 0 0 $X=3970 $Y=-5470
X33 8 M1_PO_CDNS_7654617506820 $T=4540 -5740 0 0 $X=4300 $Y=-5840
X34 5 M1_PO_CDNS_7654617506820 $T=4960 -4960 0 0 $X=4720 $Y=-5060
X35 5 M1_PO_CDNS_7654617506820 $T=4960 -2500 0 0 $X=4720 $Y=-2600
X36 1 5 9 2 6 pmos1v_CDNS_765461750688 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 2 7 3 nmos1v_CDNS_765461750689 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 9 6 7 2 pmos1v_CDNS_7654617506810 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 6 8 11 2 pmos1v_CDNS_7654617506811 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 3 7 11 2 6 pmos1v_CDNS_7654617506812 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X41 2 3 8 2 nmos1v_CDNS_7654617506813 $T=1570 -6390 0 270 $X=1370 $Y=-6840
X42 10 1 8 2 nmos1v_CDNS_7654617506813 $T=1570 -4430 0 270 $X=1370 $Y=-4880
X43 10 7 2 nmos1v_CDNS_7654617506814 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 4 1 12 2 nmos1v_CDNS_7654617506815 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 2 5 12 nmos1v_CDNS_7654617506816 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 9 8 6 2 pmos1v_CDNS_7654617506817 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 9 4 1 2 6 pmos1v_CDNS_7654617506818 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 2 8 3 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 10 8 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M2 6 4 8 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=5520 $Y=-3590 $dt=1
M3 6 5 7 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5520 $Y=-2660 $dt=1
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7654617506821                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7654617506821 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7654617506821

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7654617506822                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7654617506822 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7654617506822

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7654617506823                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7654617506823 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7654617506823

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7654617506824                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7654617506824 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7654617506824

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7654617506825                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7654617506825 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7654617506825

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7654617506826                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7654617506826 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7654617506826

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7654617506827                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7654617506827 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7654617506827

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7654617506829                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7654617506829 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7654617506829

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7654617506830                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7654617506830 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7654617506830

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7654617506831                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7654617506831 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7654617506831

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7654617506832                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7654617506832 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7654617506832

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7654617506833                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7654617506833 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7654617506833

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7654617506834                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7654617506834 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7654617506834

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506819                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506819 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 4 3 1 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506820                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506820 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39
*.DEVICECLIMB
** N=39 EP=39 FDC=54
X0 2 M4_M3_CDNS_765461750680 $T=610 4030 0 0 $X=530 $Y=3780
X1 1 M4_M3_CDNS_765461750680 $T=930 5440 0 0 $X=850 $Y=5190
X2 2 M4_M3_CDNS_765461750680 $T=2790 4030 0 0 $X=2710 $Y=3780
X3 1 M4_M3_CDNS_765461750680 $T=5580 5440 0 0 $X=5500 $Y=5190
X4 2 M4_M3_CDNS_765461750680 $T=7440 4030 0 0 $X=7360 $Y=3780
X5 10 M4_M3_CDNS_765461750680 $T=8700 3090 0 0 $X=8620 $Y=2840
X6 9 M4_M3_CDNS_765461750680 $T=10230 6380 0 0 $X=10150 $Y=6130
X7 1 M4_M3_CDNS_765461750680 $T=12090 5440 0 0 $X=12010 $Y=5190
X8 2 M4_M3_CDNS_765461750680 $T=13950 4030 0 0 $X=13870 $Y=3780
X9 10 M4_M3_CDNS_765461750680 $T=15810 3090 0 0 $X=15730 $Y=2840
X10 9 M4_M3_CDNS_765461750680 $T=18600 6380 0 0 $X=18520 $Y=6130
X11 1 M4_M3_CDNS_765461750680 $T=20460 5440 0 0 $X=20380 $Y=5190
X12 2 M4_M3_CDNS_765461750680 $T=22320 4030 0 0 $X=22240 $Y=3780
X13 10 M4_M3_CDNS_765461750680 $T=24180 3090 0 0 $X=24100 $Y=2840
X14 16 M5_M4_CDNS_765461750684 $T=3580 4500 0 0 $X=3360 $Y=4250
X15 17 M5_M4_CDNS_765461750684 $T=9160 4500 0 0 $X=8940 $Y=4250
X16 18 M5_M4_CDNS_765461750684 $T=16600 4500 0 0 $X=16380 $Y=4250
X17 19 M5_M4_CDNS_765461750684 $T=25900 4500 0 0 $X=25680 $Y=4250
X18 2 M3_M2_CDNS_765461750685 $T=610 4030 0 0 $X=530 $Y=3780
X19 1 M3_M2_CDNS_765461750685 $T=930 5440 0 0 $X=850 $Y=5190
X20 2 M3_M2_CDNS_765461750685 $T=2790 4030 0 0 $X=2710 $Y=3780
X21 7 M3_M2_CDNS_765461750685 $T=3110 3560 0 0 $X=3030 $Y=3310
X22 8 M3_M2_CDNS_765461750685 $T=4110 1490 0 0 $X=4030 $Y=1240
X23 1 M3_M2_CDNS_765461750685 $T=5580 5440 0 0 $X=5500 $Y=5190
X24 2 M3_M2_CDNS_765461750685 $T=7440 4030 0 0 $X=7360 $Y=3780
X25 10 M3_M2_CDNS_765461750685 $T=8700 3090 0 0 $X=8620 $Y=2840
X26 11 M3_M2_CDNS_765461750685 $T=9690 1490 0 0 $X=9610 $Y=1240
X27 9 M3_M2_CDNS_765461750685 $T=10230 6380 0 0 $X=10150 $Y=6130
X28 1 M3_M2_CDNS_765461750685 $T=12090 5440 0 0 $X=12010 $Y=5190
X29 2 M3_M2_CDNS_765461750685 $T=13950 4030 0 0 $X=13870 $Y=3780
X30 10 M3_M2_CDNS_765461750685 $T=15810 3090 0 0 $X=15730 $Y=2840
X31 13 M3_M2_CDNS_765461750685 $T=17130 1490 0 0 $X=17050 $Y=1240
X32 14 M3_M2_CDNS_765461750685 $T=17490 2630 0 0 $X=17410 $Y=2380
X33 9 M3_M2_CDNS_765461750685 $T=18600 6380 0 0 $X=18520 $Y=6130
X34 1 M3_M2_CDNS_765461750685 $T=20460 5440 0 0 $X=20380 $Y=5190
X35 2 M3_M2_CDNS_765461750685 $T=22320 4030 0 0 $X=22240 $Y=3780
X36 10 M3_M2_CDNS_765461750685 $T=24180 3090 0 0 $X=24100 $Y=2840
X37 15 M3_M2_CDNS_765461750685 $T=26430 1490 0 0 $X=26350 $Y=1240
X38 16 M4_M3_CDNS_765461750686 $T=3580 4500 0 0 $X=3360 $Y=4250
X39 17 M4_M3_CDNS_765461750686 $T=9160 4500 0 0 $X=8940 $Y=4250
X40 18 M4_M3_CDNS_765461750686 $T=16600 4500 0 0 $X=16380 $Y=4250
X41 19 M4_M3_CDNS_765461750686 $T=25900 4500 0 0 $X=25680 $Y=4250
X42 16 M3_M2_CDNS_765461750687 $T=3580 4500 0 0 $X=3360 $Y=4250
X43 17 M3_M2_CDNS_765461750687 $T=9160 4500 0 0 $X=8940 $Y=4250
X44 18 M3_M2_CDNS_765461750687 $T=16600 4500 0 0 $X=16380 $Y=4250
X45 19 M3_M2_CDNS_765461750687 $T=25900 4500 0 0 $X=25680 $Y=4250
X46 16 M2_M1_CDNS_765461750688 $T=3580 4500 0 0 $X=3360 $Y=4250
X47 17 M2_M1_CDNS_765461750688 $T=9160 4500 0 0 $X=8940 $Y=4250
X48 18 M2_M1_CDNS_765461750688 $T=16600 4500 0 0 $X=16380 $Y=4250
X49 19 M2_M1_CDNS_765461750688 $T=25900 4500 0 0 $X=25680 $Y=4250
X50 7 M4_M3_CDNS_7654617506811 $T=3110 3560 0 0 $X=3030 $Y=3310
X51 8 M4_M3_CDNS_7654617506811 $T=4110 1490 0 0 $X=4030 $Y=1240
X52 11 M4_M3_CDNS_7654617506811 $T=9690 1490 0 0 $X=9610 $Y=1240
X53 13 M4_M3_CDNS_7654617506811 $T=17130 1490 0 0 $X=17050 $Y=1240
X54 14 M4_M3_CDNS_7654617506811 $T=17490 2630 0 0 $X=17410 $Y=2380
X55 15 M4_M3_CDNS_7654617506811 $T=26430 1490 0 0 $X=26350 $Y=1240
X56 3 M3_M2_CDNS_7654617506813 $T=250 4970 0 90 $X=0 $Y=4890
X57 3 M3_M2_CDNS_7654617506813 $T=1860 4970 0 0 $X=1780 $Y=4720
X58 6 M3_M2_CDNS_7654617506813 $T=4650 5910 0 0 $X=4570 $Y=5660
X59 3 M3_M2_CDNS_7654617506813 $T=6510 4970 0 0 $X=6430 $Y=4720
X60 7 M3_M2_CDNS_7654617506813 $T=8370 3560 0 0 $X=8290 $Y=3310
X61 6 M3_M2_CDNS_7654617506813 $T=11160 5910 0 0 $X=11080 $Y=5660
X62 3 M3_M2_CDNS_7654617506813 $T=13020 4970 0 0 $X=12940 $Y=4720
X63 7 M3_M2_CDNS_7654617506813 $T=14880 3560 0 0 $X=14800 $Y=3310
X64 12 M3_M2_CDNS_7654617506813 $T=17670 6850 0 0 $X=17590 $Y=6600
X65 6 M3_M2_CDNS_7654617506813 $T=19530 5910 0 0 $X=19450 $Y=5660
X66 3 M3_M2_CDNS_7654617506813 $T=21390 4970 0 0 $X=21310 $Y=4720
X67 7 M3_M2_CDNS_7654617506813 $T=23250 3560 0 0 $X=23170 $Y=3310
X68 14 M3_M2_CDNS_7654617506813 $T=25110 2620 0 0 $X=25030 $Y=2370
X69 3 M2_M1_CDNS_7654617506814 $T=250 4970 0 90 $X=0 $Y=4890
X70 4 4 2 20 5 pmos1v_CDNS_765461750686 $T=2980 8370 1 180 $X=2470 $Y=8170
X71 4 4 16 8 5 pmos1v_CDNS_765461750686 $T=3820 8370 0 0 $X=3400 $Y=8170
X72 4 4 6 17 5 pmos1v_CDNS_765461750686 $T=4750 8370 0 0 $X=4330 $Y=8170
X73 21 4 3 17 5 pmos1v_CDNS_765461750686 $T=6700 8370 1 180 $X=6190 $Y=8170
X74 22 4 2 21 5 pmos1v_CDNS_765461750686 $T=7630 8370 1 180 $X=7120 $Y=8170
X75 4 4 7 22 5 pmos1v_CDNS_765461750686 $T=8560 8370 1 180 $X=8050 $Y=8170
X76 4 4 17 11 5 pmos1v_CDNS_765461750686 $T=9400 8370 0 0 $X=8980 $Y=8170
X77 4 4 9 18 5 pmos1v_CDNS_765461750686 $T=10330 8370 0 0 $X=9910 $Y=8170
X78 23 4 6 18 5 pmos1v_CDNS_765461750686 $T=11350 8370 1 180 $X=10840 $Y=8170
X79 24 4 1 18 5 pmos1v_CDNS_765461750686 $T=12280 8370 1 180 $X=11770 $Y=8170
X80 25 4 3 18 5 pmos1v_CDNS_765461750686 $T=13210 8370 1 180 $X=12700 $Y=8170
X81 24 4 2 25 5 pmos1v_CDNS_765461750686 $T=14140 8370 1 180 $X=13630 $Y=8170
X82 23 4 7 24 5 pmos1v_CDNS_765461750686 $T=15070 8370 1 180 $X=14560 $Y=8170
X83 4 4 10 23 5 pmos1v_CDNS_765461750686 $T=16000 8370 1 180 $X=15490 $Y=8170
X84 4 4 12 19 5 pmos1v_CDNS_765461750686 $T=17770 8370 0 0 $X=17350 $Y=8170
X85 26 4 6 19 5 pmos1v_CDNS_765461750686 $T=19720 8370 1 180 $X=19210 $Y=8170
X86 27 4 1 19 5 pmos1v_CDNS_765461750686 $T=20650 8370 1 180 $X=20140 $Y=8170
X87 27 4 2 28 5 pmos1v_CDNS_765461750686 $T=22510 8370 1 180 $X=22000 $Y=8170
X88 26 4 7 27 5 pmos1v_CDNS_765461750686 $T=23440 8370 1 180 $X=22930 $Y=8170
X89 4 4 14 29 5 pmos1v_CDNS_765461750686 $T=25300 8370 1 180 $X=24790 $Y=8170
X90 4 4 19 15 5 pmos1v_CDNS_765461750686 $T=26140 8370 0 0 $X=25720 $Y=8170
X91 5 5 1 30 nmos1v_CDNS_765461750687 $T=1030 800 0 0 $X=610 $Y=240
X92 30 5 3 16 nmos1v_CDNS_765461750687 $T=1960 800 0 0 $X=1540 $Y=240
X93 5 5 6 31 nmos1v_CDNS_765461750687 $T=4750 800 0 0 $X=4330 $Y=240
X94 31 5 2 17 nmos1v_CDNS_765461750687 $T=7540 800 0 0 $X=7120 $Y=240
X95 5 5 7 17 nmos1v_CDNS_765461750687 $T=8560 800 1 180 $X=8050 $Y=240
X96 5 5 17 11 nmos1v_CDNS_765461750687 $T=9400 800 0 0 $X=8980 $Y=240
X97 32 5 1 33 nmos1v_CDNS_765461750687 $T=12190 800 0 0 $X=11770 $Y=240
X98 33 5 3 18 nmos1v_CDNS_765461750687 $T=13120 800 0 0 $X=12700 $Y=240
X99 34 5 7 18 nmos1v_CDNS_765461750687 $T=14980 800 0 0 $X=14560 $Y=240
X100 5 5 10 18 nmos1v_CDNS_765461750687 $T=16000 800 1 180 $X=15490 $Y=240
X101 5 5 18 13 nmos1v_CDNS_765461750687 $T=16840 800 0 0 $X=16420 $Y=240
X102 35 5 9 36 nmos1v_CDNS_765461750687 $T=18700 800 0 0 $X=18280 $Y=240
X103 36 5 7 19 nmos1v_CDNS_765461750687 $T=23350 800 0 0 $X=22930 $Y=240
X104 5 5 19 15 nmos1v_CDNS_765461750687 $T=26140 800 0 0 $X=25720 $Y=240
X105 1 M4_M3_CDNS_7654617506821 $T=80 5580 0 0 $X=0 $Y=5190
X106 16 M4_M3_CDNS_7654617506821 $T=1540 7840 0 0 $X=1460 $Y=7450
X107 6 M4_M3_CDNS_7654617506821 $T=2130 6050 0 0 $X=2050 $Y=5660
X108 16 M4_M3_CDNS_7654617506821 $T=2470 1570 0 0 $X=2390 $Y=1180
X109 17 M4_M3_CDNS_7654617506821 $T=5260 7840 0 0 $X=5180 $Y=7450
X110 17 M4_M3_CDNS_7654617506821 $T=6450 7840 0 0 $X=6370 $Y=7450
X111 17 M4_M3_CDNS_7654617506821 $T=6860 1570 0 0 $X=6780 $Y=1180
X112 9 M4_M3_CDNS_7654617506821 $T=7710 6520 0 0 $X=7630 $Y=6130
X113 17 M4_M3_CDNS_7654617506821 $T=8050 1570 0 0 $X=7970 $Y=1180
X114 18 M4_M3_CDNS_7654617506821 $T=10840 7840 0 0 $X=10760 $Y=7450
X115 18 M4_M3_CDNS_7654617506821 $T=12030 7840 0 0 $X=11950 $Y=7450
X116 18 M4_M3_CDNS_7654617506821 $T=12960 7840 0 0 $X=12880 $Y=7450
X117 18 M4_M3_CDNS_7654617506821 $T=13370 1570 0 0 $X=13290 $Y=1180
X118 18 M4_M3_CDNS_7654617506821 $T=14300 1570 0 0 $X=14220 $Y=1180
X119 18 M4_M3_CDNS_7654617506821 $T=15490 1570 0 0 $X=15410 $Y=1180
X120 12 M4_M3_CDNS_7654617506821 $T=16080 6990 0 0 $X=16000 $Y=6600
X121 19 M4_M3_CDNS_7654617506821 $T=18280 7840 0 0 $X=18200 $Y=7450
X122 19 M4_M3_CDNS_7654617506821 $T=19470 7840 0 0 $X=19390 $Y=7450
X123 19 M4_M3_CDNS_7654617506821 $T=20400 7840 0 0 $X=20320 $Y=7450
X124 19 M4_M3_CDNS_7654617506821 $T=21330 7840 0 0 $X=21250 $Y=7450
X125 19 M4_M3_CDNS_7654617506821 $T=21740 1570 0 0 $X=21660 $Y=1180
X126 19 M4_M3_CDNS_7654617506821 $T=22670 1570 0 0 $X=22590 $Y=1180
X127 19 M4_M3_CDNS_7654617506821 $T=23600 1570 0 0 $X=23520 $Y=1180
X128 19 M4_M3_CDNS_7654617506821 $T=24790 1570 0 0 $X=24710 $Y=1180
X129 16 M7_M6_CDNS_7654617506822 $T=1540 7840 0 0 $X=1460 $Y=7450
X130 16 M7_M6_CDNS_7654617506822 $T=2470 1570 0 0 $X=2390 $Y=1180
X131 17 M7_M6_CDNS_7654617506822 $T=5260 7840 0 0 $X=5180 $Y=7450
X132 17 M7_M6_CDNS_7654617506822 $T=6450 7840 0 0 $X=6370 $Y=7450
X133 17 M7_M6_CDNS_7654617506822 $T=6860 1570 0 0 $X=6780 $Y=1180
X134 17 M7_M6_CDNS_7654617506822 $T=8050 1570 0 0 $X=7970 $Y=1180
X135 18 M7_M6_CDNS_7654617506822 $T=10840 7840 0 0 $X=10760 $Y=7450
X136 18 M7_M6_CDNS_7654617506822 $T=12030 7840 0 0 $X=11950 $Y=7450
X137 18 M7_M6_CDNS_7654617506822 $T=12960 7840 0 0 $X=12880 $Y=7450
X138 18 M7_M6_CDNS_7654617506822 $T=13370 1570 0 0 $X=13290 $Y=1180
X139 18 M7_M6_CDNS_7654617506822 $T=14300 1570 0 0 $X=14220 $Y=1180
X140 18 M7_M6_CDNS_7654617506822 $T=15490 1570 0 0 $X=15410 $Y=1180
X141 19 M7_M6_CDNS_7654617506822 $T=18280 7840 0 0 $X=18200 $Y=7450
X142 19 M7_M6_CDNS_7654617506822 $T=19470 7840 0 0 $X=19390 $Y=7450
X143 19 M7_M6_CDNS_7654617506822 $T=20400 7840 0 0 $X=20320 $Y=7450
X144 19 M7_M6_CDNS_7654617506822 $T=21330 7840 0 0 $X=21250 $Y=7450
X145 19 M7_M6_CDNS_7654617506822 $T=21740 1570 0 0 $X=21660 $Y=1180
X146 19 M7_M6_CDNS_7654617506822 $T=22670 1570 0 0 $X=22590 $Y=1180
X147 19 M7_M6_CDNS_7654617506822 $T=23600 1570 0 0 $X=23520 $Y=1180
X148 19 M7_M6_CDNS_7654617506822 $T=24790 1570 0 0 $X=24710 $Y=1180
X149 16 M1_PO_CDNS_7654617506823 $T=3580 4500 0 0 $X=3340 $Y=4250
X150 17 M1_PO_CDNS_7654617506823 $T=9160 4500 0 0 $X=8920 $Y=4250
X151 18 M1_PO_CDNS_7654617506823 $T=16600 4500 0 0 $X=16360 $Y=4250
X152 16 M6_M5_CDNS_7654617506824 $T=3580 4500 0 0 $X=3360 $Y=4250
X153 17 M6_M5_CDNS_7654617506824 $T=9160 4500 0 0 $X=8940 $Y=4250
X154 18 M6_M5_CDNS_7654617506824 $T=16600 4500 0 0 $X=16380 $Y=4250
X155 19 M6_M5_CDNS_7654617506824 $T=25900 4500 0 0 $X=25680 $Y=4250
X156 2 M5_M4_CDNS_7654617506825 $T=610 4030 0 0 $X=530 $Y=3780
X157 1 M5_M4_CDNS_7654617506825 $T=930 5440 0 0 $X=850 $Y=5190
X158 2 M5_M4_CDNS_7654617506825 $T=2790 4030 0 0 $X=2710 $Y=3780
X159 1 M5_M4_CDNS_7654617506825 $T=5580 5440 0 0 $X=5500 $Y=5190
X160 2 M5_M4_CDNS_7654617506825 $T=7440 4030 0 0 $X=7360 $Y=3780
X161 10 M5_M4_CDNS_7654617506825 $T=8700 3090 0 0 $X=8620 $Y=2840
X162 9 M5_M4_CDNS_7654617506825 $T=10230 6380 0 0 $X=10150 $Y=6130
X163 1 M5_M4_CDNS_7654617506825 $T=12090 5440 0 0 $X=12010 $Y=5190
X164 2 M5_M4_CDNS_7654617506825 $T=13950 4030 0 0 $X=13870 $Y=3780
X165 10 M5_M4_CDNS_7654617506825 $T=15810 3090 0 0 $X=15730 $Y=2840
X166 9 M5_M4_CDNS_7654617506825 $T=18600 6380 0 0 $X=18520 $Y=6130
X167 1 M5_M4_CDNS_7654617506825 $T=20460 5440 0 0 $X=20380 $Y=5190
X168 2 M5_M4_CDNS_7654617506825 $T=22320 4030 0 0 $X=22240 $Y=3780
X169 10 M5_M4_CDNS_7654617506825 $T=24180 3090 0 0 $X=24100 $Y=2840
X170 1 M1_PO_CDNS_7654617506826 $T=930 5440 0 0 $X=830 $Y=5190
X171 3 M1_PO_CDNS_7654617506826 $T=1860 4970 0 0 $X=1760 $Y=4720
X172 2 M1_PO_CDNS_7654617506826 $T=2790 4030 0 0 $X=2690 $Y=3780
X173 6 M1_PO_CDNS_7654617506826 $T=4650 5910 0 0 $X=4550 $Y=5660
X174 1 M1_PO_CDNS_7654617506826 $T=5580 5440 0 0 $X=5480 $Y=5190
X175 3 M1_PO_CDNS_7654617506826 $T=6510 4970 0 0 $X=6410 $Y=4720
X176 2 M1_PO_CDNS_7654617506826 $T=7440 4030 0 0 $X=7340 $Y=3780
X177 7 M1_PO_CDNS_7654617506826 $T=8370 3560 0 0 $X=8270 $Y=3310
X178 9 M1_PO_CDNS_7654617506826 $T=10230 6380 0 0 $X=10130 $Y=6130
X179 6 M1_PO_CDNS_7654617506826 $T=11160 5910 0 0 $X=11060 $Y=5660
X180 1 M1_PO_CDNS_7654617506826 $T=12090 5440 0 0 $X=11990 $Y=5190
X181 3 M1_PO_CDNS_7654617506826 $T=13020 4970 0 0 $X=12920 $Y=4720
X182 2 M1_PO_CDNS_7654617506826 $T=13950 4030 0 0 $X=13850 $Y=3780
X183 7 M1_PO_CDNS_7654617506826 $T=14880 3560 0 0 $X=14780 $Y=3310
X184 10 M1_PO_CDNS_7654617506826 $T=15810 3090 0 0 $X=15710 $Y=2840
X185 12 M1_PO_CDNS_7654617506826 $T=17670 6850 0 0 $X=17570 $Y=6600
X186 9 M1_PO_CDNS_7654617506826 $T=18600 6380 0 0 $X=18500 $Y=6130
X187 6 M1_PO_CDNS_7654617506826 $T=19530 5910 0 0 $X=19430 $Y=5660
X188 1 M1_PO_CDNS_7654617506826 $T=20460 5440 0 0 $X=20360 $Y=5190
X189 3 M1_PO_CDNS_7654617506826 $T=21390 4970 0 0 $X=21290 $Y=4720
X190 2 M1_PO_CDNS_7654617506826 $T=22320 4030 0 0 $X=22220 $Y=3780
X191 7 M1_PO_CDNS_7654617506826 $T=23250 3560 0 0 $X=23150 $Y=3310
X192 10 M1_PO_CDNS_7654617506826 $T=24180 3090 0 0 $X=24080 $Y=2840
X193 14 M1_PO_CDNS_7654617506826 $T=25110 2620 0 0 $X=25010 $Y=2370
X194 2 M2_M1_CDNS_7654617506827 $T=610 4030 0 0 $X=530 $Y=3780
X195 1 M2_M1_CDNS_7654617506827 $T=930 5440 0 0 $X=850 $Y=5190
X196 3 M2_M1_CDNS_7654617506827 $T=1860 4970 0 0 $X=1780 $Y=4720
X197 2 M2_M1_CDNS_7654617506827 $T=2790 4030 0 0 $X=2710 $Y=3780
X198 7 M2_M1_CDNS_7654617506827 $T=3110 3560 0 0 $X=3030 $Y=3310
X199 8 M2_M1_CDNS_7654617506827 $T=4110 1490 0 0 $X=4030 $Y=1240
X200 6 M2_M1_CDNS_7654617506827 $T=4650 5910 0 0 $X=4570 $Y=5660
X201 1 M2_M1_CDNS_7654617506827 $T=5580 5440 0 0 $X=5500 $Y=5190
X202 3 M2_M1_CDNS_7654617506827 $T=6510 4970 0 0 $X=6430 $Y=4720
X203 2 M2_M1_CDNS_7654617506827 $T=7440 4030 0 0 $X=7360 $Y=3780
X204 7 M2_M1_CDNS_7654617506827 $T=8370 3560 0 0 $X=8290 $Y=3310
X205 10 M2_M1_CDNS_7654617506827 $T=8700 3090 0 0 $X=8620 $Y=2840
X206 11 M2_M1_CDNS_7654617506827 $T=9690 1490 0 0 $X=9610 $Y=1240
X207 9 M2_M1_CDNS_7654617506827 $T=10230 6380 0 0 $X=10150 $Y=6130
X208 6 M2_M1_CDNS_7654617506827 $T=11160 5910 0 0 $X=11080 $Y=5660
X209 1 M2_M1_CDNS_7654617506827 $T=12090 5440 0 0 $X=12010 $Y=5190
X210 3 M2_M1_CDNS_7654617506827 $T=13020 4970 0 0 $X=12940 $Y=4720
X211 2 M2_M1_CDNS_7654617506827 $T=13950 4030 0 0 $X=13870 $Y=3780
X212 7 M2_M1_CDNS_7654617506827 $T=14880 3560 0 0 $X=14800 $Y=3310
X213 10 M2_M1_CDNS_7654617506827 $T=15810 3090 0 0 $X=15730 $Y=2840
X214 13 M2_M1_CDNS_7654617506827 $T=17130 1490 0 0 $X=17050 $Y=1240
X215 14 M2_M1_CDNS_7654617506827 $T=17490 2630 0 0 $X=17410 $Y=2380
X216 12 M2_M1_CDNS_7654617506827 $T=17670 6850 0 0 $X=17590 $Y=6600
X217 9 M2_M1_CDNS_7654617506827 $T=18600 6380 0 0 $X=18520 $Y=6130
X218 6 M2_M1_CDNS_7654617506827 $T=19530 5910 0 0 $X=19450 $Y=5660
X219 1 M2_M1_CDNS_7654617506827 $T=20460 5440 0 0 $X=20380 $Y=5190
X220 3 M2_M1_CDNS_7654617506827 $T=21390 4970 0 0 $X=21310 $Y=4720
X221 2 M2_M1_CDNS_7654617506827 $T=22320 4030 0 0 $X=22240 $Y=3780
X222 7 M2_M1_CDNS_7654617506827 $T=23250 3560 0 0 $X=23170 $Y=3310
X223 10 M2_M1_CDNS_7654617506827 $T=24180 3090 0 0 $X=24100 $Y=2840
X224 14 M2_M1_CDNS_7654617506827 $T=25110 2620 0 0 $X=25030 $Y=2370
X225 15 M2_M1_CDNS_7654617506827 $T=26430 1490 0 0 $X=26350 $Y=1240
X226 1 M2_M1_CDNS_7654617506829 $T=80 5580 0 0 $X=0 $Y=5190
X227 16 M2_M1_CDNS_7654617506829 $T=1540 7840 0 0 $X=1460 $Y=7450
X228 6 M2_M1_CDNS_7654617506829 $T=2130 6050 0 0 $X=2050 $Y=5660
X229 16 M2_M1_CDNS_7654617506829 $T=2470 1570 0 0 $X=2390 $Y=1180
X230 17 M2_M1_CDNS_7654617506829 $T=5260 7840 0 0 $X=5180 $Y=7450
X231 17 M2_M1_CDNS_7654617506829 $T=6450 7840 0 0 $X=6370 $Y=7450
X232 17 M2_M1_CDNS_7654617506829 $T=6860 1570 0 0 $X=6780 $Y=1180
X233 9 M2_M1_CDNS_7654617506829 $T=7710 6520 0 0 $X=7630 $Y=6130
X234 17 M2_M1_CDNS_7654617506829 $T=8050 1570 0 0 $X=7970 $Y=1180
X235 18 M2_M1_CDNS_7654617506829 $T=10840 7840 0 0 $X=10760 $Y=7450
X236 18 M2_M1_CDNS_7654617506829 $T=12030 7840 0 0 $X=11950 $Y=7450
X237 18 M2_M1_CDNS_7654617506829 $T=12960 7840 0 0 $X=12880 $Y=7450
X238 18 M2_M1_CDNS_7654617506829 $T=13370 1570 0 0 $X=13290 $Y=1180
X239 18 M2_M1_CDNS_7654617506829 $T=14300 1570 0 0 $X=14220 $Y=1180
X240 18 M2_M1_CDNS_7654617506829 $T=15490 1570 0 0 $X=15410 $Y=1180
X241 12 M2_M1_CDNS_7654617506829 $T=16080 6990 0 0 $X=16000 $Y=6600
X242 19 M2_M1_CDNS_7654617506829 $T=18280 7840 0 0 $X=18200 $Y=7450
X243 19 M2_M1_CDNS_7654617506829 $T=19470 7840 0 0 $X=19390 $Y=7450
X244 19 M2_M1_CDNS_7654617506829 $T=20400 7840 0 0 $X=20320 $Y=7450
X245 19 M2_M1_CDNS_7654617506829 $T=21330 7840 0 0 $X=21250 $Y=7450
X246 19 M2_M1_CDNS_7654617506829 $T=21740 1570 0 0 $X=21660 $Y=1180
X247 19 M2_M1_CDNS_7654617506829 $T=22670 1570 0 0 $X=22590 $Y=1180
X248 19 M2_M1_CDNS_7654617506829 $T=23600 1570 0 0 $X=23520 $Y=1180
X249 19 M2_M1_CDNS_7654617506829 $T=24790 1570 0 0 $X=24710 $Y=1180
X250 16 M7_M6_CDNS_7654617506830 $T=3580 4500 0 0 $X=3360 $Y=4250
X251 17 M7_M6_CDNS_7654617506830 $T=9160 4500 0 0 $X=8940 $Y=4250
X252 18 M7_M6_CDNS_7654617506830 $T=16600 4500 0 0 $X=16380 $Y=4250
X253 19 M7_M6_CDNS_7654617506830 $T=25900 4500 0 0 $X=25680 $Y=4250
X254 16 M6_M5_CDNS_7654617506831 $T=1540 7840 0 0 $X=1460 $Y=7450
X255 16 M6_M5_CDNS_7654617506831 $T=2470 1570 0 0 $X=2390 $Y=1180
X256 17 M6_M5_CDNS_7654617506831 $T=5260 7840 0 0 $X=5180 $Y=7450
X257 17 M6_M5_CDNS_7654617506831 $T=6450 7840 0 0 $X=6370 $Y=7450
X258 17 M6_M5_CDNS_7654617506831 $T=6860 1570 0 0 $X=6780 $Y=1180
X259 17 M6_M5_CDNS_7654617506831 $T=8050 1570 0 0 $X=7970 $Y=1180
X260 18 M6_M5_CDNS_7654617506831 $T=10840 7840 0 0 $X=10760 $Y=7450
X261 18 M6_M5_CDNS_7654617506831 $T=12030 7840 0 0 $X=11950 $Y=7450
X262 18 M6_M5_CDNS_7654617506831 $T=12960 7840 0 0 $X=12880 $Y=7450
X263 18 M6_M5_CDNS_7654617506831 $T=13370 1570 0 0 $X=13290 $Y=1180
X264 18 M6_M5_CDNS_7654617506831 $T=14300 1570 0 0 $X=14220 $Y=1180
X265 18 M6_M5_CDNS_7654617506831 $T=15490 1570 0 0 $X=15410 $Y=1180
X266 19 M6_M5_CDNS_7654617506831 $T=18280 7840 0 0 $X=18200 $Y=7450
X267 19 M6_M5_CDNS_7654617506831 $T=19470 7840 0 0 $X=19390 $Y=7450
X268 19 M6_M5_CDNS_7654617506831 $T=20400 7840 0 0 $X=20320 $Y=7450
X269 19 M6_M5_CDNS_7654617506831 $T=21330 7840 0 0 $X=21250 $Y=7450
X270 19 M6_M5_CDNS_7654617506831 $T=21740 1570 0 0 $X=21660 $Y=1180
X271 19 M6_M5_CDNS_7654617506831 $T=22670 1570 0 0 $X=22590 $Y=1180
X272 19 M6_M5_CDNS_7654617506831 $T=23600 1570 0 0 $X=23520 $Y=1180
X273 19 M6_M5_CDNS_7654617506831 $T=24790 1570 0 0 $X=24710 $Y=1180
X274 1 M6_M5_CDNS_7654617506832 $T=80 5580 0 0 $X=0 $Y=5190
X275 6 M6_M5_CDNS_7654617506832 $T=2130 6050 0 0 $X=2050 $Y=5660
X276 9 M6_M5_CDNS_7654617506832 $T=7710 6520 0 0 $X=7630 $Y=6130
X277 12 M6_M5_CDNS_7654617506832 $T=16080 6990 0 0 $X=16000 $Y=6600
X278 1 M3_M2_CDNS_7654617506833 $T=80 5580 0 0 $X=0 $Y=5190
X279 16 M3_M2_CDNS_7654617506833 $T=1540 7840 0 0 $X=1460 $Y=7450
X280 6 M3_M2_CDNS_7654617506833 $T=2130 6050 0 0 $X=2050 $Y=5660
X281 16 M3_M2_CDNS_7654617506833 $T=2470 1570 0 0 $X=2390 $Y=1180
X282 17 M3_M2_CDNS_7654617506833 $T=5260 7840 0 0 $X=5180 $Y=7450
X283 17 M3_M2_CDNS_7654617506833 $T=6450 7840 0 0 $X=6370 $Y=7450
X284 17 M3_M2_CDNS_7654617506833 $T=6860 1570 0 0 $X=6780 $Y=1180
X285 9 M3_M2_CDNS_7654617506833 $T=7710 6520 0 0 $X=7630 $Y=6130
X286 17 M3_M2_CDNS_7654617506833 $T=8050 1570 0 0 $X=7970 $Y=1180
X287 18 M3_M2_CDNS_7654617506833 $T=10840 7840 0 0 $X=10760 $Y=7450
X288 18 M3_M2_CDNS_7654617506833 $T=12030 7840 0 0 $X=11950 $Y=7450
X289 18 M3_M2_CDNS_7654617506833 $T=12960 7840 0 0 $X=12880 $Y=7450
X290 18 M3_M2_CDNS_7654617506833 $T=13370 1570 0 0 $X=13290 $Y=1180
X291 18 M3_M2_CDNS_7654617506833 $T=14300 1570 0 0 $X=14220 $Y=1180
X292 18 M3_M2_CDNS_7654617506833 $T=15490 1570 0 0 $X=15410 $Y=1180
X293 12 M3_M2_CDNS_7654617506833 $T=16080 6990 0 0 $X=16000 $Y=6600
X294 19 M3_M2_CDNS_7654617506833 $T=18280 7840 0 0 $X=18200 $Y=7450
X295 19 M3_M2_CDNS_7654617506833 $T=19470 7840 0 0 $X=19390 $Y=7450
X296 19 M3_M2_CDNS_7654617506833 $T=20400 7840 0 0 $X=20320 $Y=7450
X297 19 M3_M2_CDNS_7654617506833 $T=21330 7840 0 0 $X=21250 $Y=7450
X298 19 M3_M2_CDNS_7654617506833 $T=21740 1570 0 0 $X=21660 $Y=1180
X299 19 M3_M2_CDNS_7654617506833 $T=22670 1570 0 0 $X=22590 $Y=1180
X300 19 M3_M2_CDNS_7654617506833 $T=23600 1570 0 0 $X=23520 $Y=1180
X301 19 M3_M2_CDNS_7654617506833 $T=24790 1570 0 0 $X=24710 $Y=1180
X302 1 M5_M4_CDNS_7654617506834 $T=80 5580 0 0 $X=0 $Y=5190
X303 16 M5_M4_CDNS_7654617506834 $T=1540 7840 0 0 $X=1460 $Y=7450
X304 6 M5_M4_CDNS_7654617506834 $T=2130 6050 0 0 $X=2050 $Y=5660
X305 16 M5_M4_CDNS_7654617506834 $T=2470 1570 0 0 $X=2390 $Y=1180
X306 17 M5_M4_CDNS_7654617506834 $T=5260 7840 0 0 $X=5180 $Y=7450
X307 17 M5_M4_CDNS_7654617506834 $T=6450 7840 0 0 $X=6370 $Y=7450
X308 17 M5_M4_CDNS_7654617506834 $T=6860 1570 0 0 $X=6780 $Y=1180
X309 9 M5_M4_CDNS_7654617506834 $T=7710 6520 0 0 $X=7630 $Y=6130
X310 17 M5_M4_CDNS_7654617506834 $T=8050 1570 0 0 $X=7970 $Y=1180
X311 18 M5_M4_CDNS_7654617506834 $T=10840 7840 0 0 $X=10760 $Y=7450
X312 18 M5_M4_CDNS_7654617506834 $T=12030 7840 0 0 $X=11950 $Y=7450
X313 18 M5_M4_CDNS_7654617506834 $T=12960 7840 0 0 $X=12880 $Y=7450
X314 18 M5_M4_CDNS_7654617506834 $T=13370 1570 0 0 $X=13290 $Y=1180
X315 18 M5_M4_CDNS_7654617506834 $T=14300 1570 0 0 $X=14220 $Y=1180
X316 18 M5_M4_CDNS_7654617506834 $T=15490 1570 0 0 $X=15410 $Y=1180
X317 12 M5_M4_CDNS_7654617506834 $T=16080 6990 0 0 $X=16000 $Y=6600
X318 19 M5_M4_CDNS_7654617506834 $T=18280 7840 0 0 $X=18200 $Y=7450
X319 19 M5_M4_CDNS_7654617506834 $T=19470 7840 0 0 $X=19390 $Y=7450
X320 19 M5_M4_CDNS_7654617506834 $T=20400 7840 0 0 $X=20320 $Y=7450
X321 19 M5_M4_CDNS_7654617506834 $T=21330 7840 0 0 $X=21250 $Y=7450
X322 19 M5_M4_CDNS_7654617506834 $T=21740 1570 0 0 $X=21660 $Y=1180
X323 19 M5_M4_CDNS_7654617506834 $T=22670 1570 0 0 $X=22590 $Y=1180
X324 19 M5_M4_CDNS_7654617506834 $T=23600 1570 0 0 $X=23520 $Y=1180
X325 19 M5_M4_CDNS_7654617506834 $T=24790 1570 0 0 $X=24710 $Y=1180
X326 4 4 1 16 5 pmos1v_CDNS_7654617506819 $T=1030 8610 1 0 $X=610 $Y=8170
X327 20 4 3 16 5 pmos1v_CDNS_7654617506819 $T=2050 8610 0 180 $X=1540 $Y=8170
X328 22 4 1 17 5 pmos1v_CDNS_7654617506819 $T=5770 8610 0 180 $X=5260 $Y=8170
X329 4 4 18 13 5 pmos1v_CDNS_7654617506819 $T=16840 8610 1 0 $X=16420 $Y=8170
X330 29 4 9 19 5 pmos1v_CDNS_7654617506819 $T=18790 8610 0 180 $X=18280 $Y=8170
X331 28 4 3 19 5 pmos1v_CDNS_7654617506819 $T=21580 8610 0 180 $X=21070 $Y=8170
X332 29 4 10 26 5 pmos1v_CDNS_7654617506819 $T=24370 8610 0 180 $X=23860 $Y=8170
X333 5 5 2 16 nmos1v_CDNS_7654617506820 $T=2980 1040 0 180 $X=2470 $Y=240
X334 5 5 16 8 nmos1v_CDNS_7654617506820 $T=3820 1040 1 0 $X=3400 $Y=240
X335 31 5 1 37 nmos1v_CDNS_7654617506820 $T=5680 1040 1 0 $X=5260 $Y=240
X336 37 5 3 17 nmos1v_CDNS_7654617506820 $T=6610 1040 1 0 $X=6190 $Y=240
X337 5 5 9 34 nmos1v_CDNS_7654617506820 $T=10330 1040 1 0 $X=9910 $Y=240
X338 34 5 6 32 nmos1v_CDNS_7654617506820 $T=11260 1040 1 0 $X=10840 $Y=240
X339 32 5 2 18 nmos1v_CDNS_7654617506820 $T=14050 1040 1 0 $X=13630 $Y=240
X340 5 5 12 35 nmos1v_CDNS_7654617506820 $T=17770 1040 1 0 $X=17350 $Y=240
X341 36 5 6 38 nmos1v_CDNS_7654617506820 $T=19630 1040 1 0 $X=19210 $Y=240
X342 38 5 1 39 nmos1v_CDNS_7654617506820 $T=20560 1040 1 0 $X=20140 $Y=240
X343 39 5 3 19 nmos1v_CDNS_7654617506820 $T=21490 1040 1 0 $X=21070 $Y=240
X344 38 5 2 19 nmos1v_CDNS_7654617506820 $T=22420 1040 1 0 $X=22000 $Y=240
X345 35 5 10 19 nmos1v_CDNS_7654617506820 $T=24280 1040 1 0 $X=23860 $Y=240
X346 5 5 14 19 nmos1v_CDNS_7654617506820 $T=25300 1040 0 180 $X=24790 $Y=240
M0 4 2 20 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M1 8 16 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M2 17 6 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M3 21 3 17 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M4 22 2 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M5 4 7 22 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M6 11 17 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M7 18 9 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M8 23 6 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M9 24 1 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M10 25 3 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M11 24 2 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M12 23 7 24 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M13 4 10 23 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M14 19 12 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M15 26 6 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M16 27 1 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M17 27 2 28 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M18 26 7 27 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceFinalAdder                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceFinalAdder 13 12 11 10 44 57 17 16 15 14
+ 39 38 37 34 45 58 43 42 41 40
+ 36 50 49 48 47 46 56 55 53 52
+ 51 35
** N=164 EP=32 FDC=320
X0 1 M4_M3_CDNS_765461750680 $T=150 2650 0 0 $X=70 $Y=2400
X1 2 M4_M3_CDNS_765461750680 $T=5940 2650 0 0 $X=5860 $Y=2400
X2 3 M4_M3_CDNS_765461750680 $T=16170 2650 0 0 $X=16090 $Y=2400
X3 4 M4_M3_CDNS_765461750680 $T=21750 2650 0 0 $X=21670 $Y=2400
X4 5 M4_M3_CDNS_765461750680 $T=26890 2650 0 0 $X=26810 $Y=2400
X5 6 M4_M3_CDNS_765461750680 $T=32670 2650 0 0 $X=32590 $Y=2400
X6 7 M4_M3_CDNS_765461750680 $T=40090 2650 0 0 $X=40010 $Y=2400
X7 8 M4_M3_CDNS_765461750680 $T=48440 2650 0 0 $X=48360 $Y=2400
X8 9 M4_M3_CDNS_765461750680 $T=53580 2650 0 0 $X=53500 $Y=2400
X9 1 M6_M5_CDNS_765461750681 $T=150 2650 0 0 $X=70 $Y=2400
X10 2 M6_M5_CDNS_765461750681 $T=5940 2650 0 0 $X=5860 $Y=2400
X11 3 M6_M5_CDNS_765461750681 $T=16170 2650 0 0 $X=16090 $Y=2400
X12 4 M6_M5_CDNS_765461750681 $T=21750 2650 0 0 $X=21670 $Y=2400
X13 5 M6_M5_CDNS_765461750681 $T=26890 2650 0 0 $X=26810 $Y=2400
X14 6 M6_M5_CDNS_765461750681 $T=32670 2650 0 0 $X=32590 $Y=2400
X15 7 M6_M5_CDNS_765461750681 $T=40090 2650 0 0 $X=40010 $Y=2400
X16 8 M6_M5_CDNS_765461750681 $T=48440 2650 0 0 $X=48360 $Y=2400
X17 9 M6_M5_CDNS_765461750681 $T=53580 2650 0 0 $X=53500 $Y=2400
X18 1 M5_M4_CDNS_765461750682 $T=150 2650 0 0 $X=70 $Y=2400
X19 2 M5_M4_CDNS_765461750682 $T=5940 2650 0 0 $X=5860 $Y=2400
X20 3 M5_M4_CDNS_765461750682 $T=16170 2650 0 0 $X=16090 $Y=2400
X21 4 M5_M4_CDNS_765461750682 $T=21750 2650 0 0 $X=21670 $Y=2400
X22 5 M5_M4_CDNS_765461750682 $T=26890 2650 0 0 $X=26810 $Y=2400
X23 6 M5_M4_CDNS_765461750682 $T=32670 2650 0 0 $X=32590 $Y=2400
X24 7 M5_M4_CDNS_765461750682 $T=40090 2650 0 0 $X=40010 $Y=2400
X25 8 M5_M4_CDNS_765461750682 $T=48440 2650 0 0 $X=48360 $Y=2400
X26 9 M5_M4_CDNS_765461750682 $T=53580 2650 0 0 $X=53500 $Y=2400
X27 10 M2_M1_CDNS_765461750683 $T=4820 20240 0 0 $X=4740 $Y=20110
X28 11 M2_M1_CDNS_765461750683 $T=13610 20240 0 0 $X=13530 $Y=20110
X29 12 M2_M1_CDNS_765461750683 $T=19200 20240 0 0 $X=19120 $Y=20110
X30 13 M2_M1_CDNS_765461750683 $T=31060 20240 0 0 $X=30980 $Y=20110
X31 14 M2_M1_CDNS_765461750683 $T=31510 20240 0 0 $X=31430 $Y=20110
X32 15 M2_M1_CDNS_765461750683 $T=40300 20240 0 0 $X=40220 $Y=20110
X33 16 M2_M1_CDNS_765461750683 $T=45890 20240 0 0 $X=45810 $Y=20110
X34 17 M2_M1_CDNS_765461750683 $T=57710 20240 0 0 $X=57630 $Y=20110
X35 18 M5_M4_CDNS_765461750684 $T=9340 19910 0 0 $X=9120 $Y=19660
X36 19 M5_M4_CDNS_765461750684 $T=18130 19910 0 0 $X=17910 $Y=19660
X37 20 M5_M4_CDNS_765461750684 $T=23720 19910 0 0 $X=23500 $Y=19660
X38 21 M5_M4_CDNS_765461750684 $T=26500 19910 0 0 $X=26280 $Y=19660
X39 22 M5_M4_CDNS_765461750684 $T=36030 19910 0 0 $X=35810 $Y=19660
X40 23 M5_M4_CDNS_765461750684 $T=44820 19910 0 0 $X=44600 $Y=19660
X41 24 M5_M4_CDNS_765461750684 $T=50410 19910 0 0 $X=50190 $Y=19660
X42 25 M5_M4_CDNS_765461750684 $T=53190 19910 0 0 $X=52970 $Y=19660
X43 1 M3_M2_CDNS_765461750685 $T=150 2650 0 0 $X=70 $Y=2400
X44 2 M3_M2_CDNS_765461750685 $T=5940 2650 0 0 $X=5860 $Y=2400
X45 3 M3_M2_CDNS_765461750685 $T=16170 2650 0 0 $X=16090 $Y=2400
X46 4 M3_M2_CDNS_765461750685 $T=21750 2650 0 0 $X=21670 $Y=2400
X47 5 M3_M2_CDNS_765461750685 $T=26890 2650 0 0 $X=26810 $Y=2400
X48 6 M3_M2_CDNS_765461750685 $T=32670 2650 0 0 $X=32590 $Y=2400
X49 7 M3_M2_CDNS_765461750685 $T=40090 2650 0 0 $X=40010 $Y=2400
X50 8 M3_M2_CDNS_765461750685 $T=48440 2650 0 0 $X=48360 $Y=2400
X51 9 M3_M2_CDNS_765461750685 $T=53580 2650 0 0 $X=53500 $Y=2400
X52 18 M4_M3_CDNS_765461750686 $T=9340 19910 0 0 $X=9120 $Y=19660
X53 19 M4_M3_CDNS_765461750686 $T=18130 19910 0 0 $X=17910 $Y=19660
X54 20 M4_M3_CDNS_765461750686 $T=23720 19910 0 0 $X=23500 $Y=19660
X55 21 M4_M3_CDNS_765461750686 $T=26500 19910 0 0 $X=26280 $Y=19660
X56 22 M4_M3_CDNS_765461750686 $T=36030 19910 0 0 $X=35810 $Y=19660
X57 23 M4_M3_CDNS_765461750686 $T=44820 19910 0 0 $X=44600 $Y=19660
X58 24 M4_M3_CDNS_765461750686 $T=50410 19910 0 0 $X=50190 $Y=19660
X59 25 M4_M3_CDNS_765461750686 $T=53190 19910 0 0 $X=52970 $Y=19660
X60 18 M3_M2_CDNS_765461750687 $T=9340 19910 0 0 $X=9120 $Y=19660
X61 19 M3_M2_CDNS_765461750687 $T=18130 19910 0 0 $X=17910 $Y=19660
X62 20 M3_M2_CDNS_765461750687 $T=23720 19910 0 0 $X=23500 $Y=19660
X63 21 M3_M2_CDNS_765461750687 $T=26500 19910 0 0 $X=26280 $Y=19660
X64 22 M3_M2_CDNS_765461750687 $T=36030 19910 0 0 $X=35810 $Y=19660
X65 23 M3_M2_CDNS_765461750687 $T=44820 19910 0 0 $X=44600 $Y=19660
X66 24 M3_M2_CDNS_765461750687 $T=50410 19910 0 0 $X=50190 $Y=19660
X67 25 M3_M2_CDNS_765461750687 $T=53190 19910 0 0 $X=52970 $Y=19660
X68 18 M2_M1_CDNS_765461750688 $T=9340 19910 0 0 $X=9120 $Y=19660
X69 19 M2_M1_CDNS_765461750688 $T=18130 19910 0 0 $X=17910 $Y=19660
X70 20 M2_M1_CDNS_765461750688 $T=23720 19910 0 0 $X=23500 $Y=19660
X71 21 M2_M1_CDNS_765461750688 $T=26500 19910 0 0 $X=26280 $Y=19660
X72 22 M2_M1_CDNS_765461750688 $T=36030 19910 0 0 $X=35810 $Y=19660
X73 23 M2_M1_CDNS_765461750688 $T=44820 19910 0 0 $X=44600 $Y=19660
X74 24 M2_M1_CDNS_765461750688 $T=50410 19910 0 0 $X=50190 $Y=19660
X75 25 M2_M1_CDNS_765461750688 $T=53190 19910 0 0 $X=52970 $Y=19660
X76 18 M6_M5_CDNS_765461750689 $T=9340 19910 0 0 $X=9120 $Y=19660
X77 19 M6_M5_CDNS_765461750689 $T=18130 19910 0 0 $X=17910 $Y=19660
X78 20 M6_M5_CDNS_765461750689 $T=23720 19910 0 0 $X=23500 $Y=19660
X79 21 M6_M5_CDNS_765461750689 $T=26500 19910 0 0 $X=26280 $Y=19660
X80 22 M6_M5_CDNS_765461750689 $T=36030 19910 0 0 $X=35810 $Y=19660
X81 23 M6_M5_CDNS_765461750689 $T=44820 19910 0 0 $X=44600 $Y=19660
X82 24 M6_M5_CDNS_765461750689 $T=50410 19910 0 0 $X=50190 $Y=19660
X83 25 M6_M5_CDNS_765461750689 $T=53190 19910 0 0 $X=52970 $Y=19660
X84 26 M3_M2_CDNS_7654617506810 $T=560 3210 0 0 $X=480 $Y=2960
X85 27 M3_M2_CDNS_7654617506810 $T=9840 3210 0 0 $X=9760 $Y=2960
X86 28 M3_M2_CDNS_7654617506810 $T=17280 3210 0 0 $X=17200 $Y=2960
X87 29 M3_M2_CDNS_7654617506810 $T=22860 3210 0 0 $X=22780 $Y=2960
X88 30 M3_M2_CDNS_7654617506810 $T=27230 3210 0 0 $X=27150 $Y=2960
X89 31 M3_M2_CDNS_7654617506810 $T=36530 3210 0 0 $X=36450 $Y=2960
X90 32 M3_M2_CDNS_7654617506810 $T=43970 3210 0 0 $X=43890 $Y=2960
X91 33 M3_M2_CDNS_7654617506810 $T=49550 3210 0 0 $X=49470 $Y=2960
X92 26 M4_M3_CDNS_7654617506811 $T=560 3210 0 0 $X=480 $Y=2960
X93 27 M4_M3_CDNS_7654617506811 $T=9840 3210 0 0 $X=9760 $Y=2960
X94 28 M4_M3_CDNS_7654617506811 $T=17280 3210 0 0 $X=17200 $Y=2960
X95 29 M4_M3_CDNS_7654617506811 $T=22860 3210 0 0 $X=22780 $Y=2960
X96 30 M4_M3_CDNS_7654617506811 $T=27230 3210 0 0 $X=27150 $Y=2960
X97 31 M4_M3_CDNS_7654617506811 $T=36530 3210 0 0 $X=36450 $Y=2960
X98 32 M4_M3_CDNS_7654617506811 $T=43970 3210 0 0 $X=43890 $Y=2960
X99 33 M4_M3_CDNS_7654617506811 $T=49550 3210 0 0 $X=49470 $Y=2960
X100 34 10 35 36 18 59 95 AND $T=3670 21910 0 0 $X=4740 $Y=18810
X101 37 11 35 36 19 60 96 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X102 38 12 35 36 20 61 97 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X103 39 13 35 36 21 62 98 AND $T=32210 21910 1 180 $X=26960 $Y=18810
X104 40 14 35 36 22 63 99 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X105 41 15 35 36 23 64 100 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X106 42 16 35 36 24 65 101 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X107 43 17 35 36 25 66 102 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X108 44 35 36 1 45 103 67 XOR $T=530 18810 1 0 $X=530 $Y=14110
X109 26 35 36 46 1 104 68 XOR $T=640 4700 1 0 $X=640 $Y=0
X110 10 35 36 2 34 105 69 XOR $T=4740 18810 1 0 $X=4740 $Y=14110
X111 27 35 36 47 2 106 70 XOR $T=9740 4700 0 180 $X=6020 $Y=0
X112 28 35 36 48 3 107 71 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X113 11 35 36 3 37 108 72 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X114 29 35 36 49 4 109 73 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X115 12 35 36 4 38 110 74 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X116 30 35 36 50 5 111 75 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X117 13 35 36 5 39 112 76 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X118 14 35 36 6 40 113 77 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X119 31 35 36 51 6 114 78 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X120 32 35 36 52 7 115 79 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X121 15 35 36 7 41 116 80 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X122 33 35 36 53 8 117 81 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X123 16 35 36 8 42 118 82 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X124 54 35 36 55 9 119 83 XOR $T=49650 4700 1 0 $X=49650 $Y=0
X125 17 35 36 9 43 120 84 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X126 56 36 54 57 58 35 86 85 143 121
+ 144 122 HAdder $T=62720 6180 1 90 $X=53760 $Y=6980
X127 5 21 30 35 36 4 20 29 3 19
+ 28 2 27 18 26 87 88 89 90 145
+ 147 146 148 149 150 152 153 154 151 123
+ 124 127 128 126 129 130 125 131 132 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X128 9 25 54 35 36 8 24 33 7 23
+ 32 6 31 22 30 91 92 93 94 155
+ 157 156 158 159 160 162 163 164 161 133
+ 134 137 138 136 139 140 135 141 142 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
M0 35 90 26 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M1 103 44 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=950 $Y=14910 $dt=1
M2 104 26 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=800 $dt=1
M3 151 18 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M4 1 45 44 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=1880 $Y=14910 $dt=1
M5 46 1 26 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=800 $dt=1
M6 103 67 1 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=2810 $Y=14910 $dt=1
M7 104 68 46 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=800 $dt=1
M8 35 45 67 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=3740 $Y=14910 $dt=1
M9 35 1 68 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=800 $dt=1
M10 105 10 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=14910 $dt=1
M11 59 10 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=20590 $dt=1
M12 35 34 59 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=20590 $dt=1
M13 2 34 10 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=14910 $dt=1
M14 70 2 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=800 $dt=1
M15 105 69 2 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=14910 $dt=1
M16 47 70 106 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=800 $dt=1
M17 35 34 69 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=14910 $dt=1
M18 27 2 47 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=800 $dt=1
M19 35 27 106 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=800 $dt=1
M20 71 3 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M21 108 11 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M22 60 11 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=20590 $dt=1
M23 35 37 60 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=20590 $dt=1
M24 48 71 107 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M25 3 37 11 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M26 28 3 48 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M27 108 72 3 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M28 35 28 107 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M29 35 37 72 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M30 73 4 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M31 110 12 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M32 61 12 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=20590 $dt=1
M33 49 73 109 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M34 35 38 61 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=20590 $dt=1
M35 4 38 12 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M36 29 4 49 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M37 110 74 4 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M38 35 29 109 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M39 35 38 74 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M40 75 5 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M41 50 75 111 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M42 30 5 50 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M43 35 30 111 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M44 35 94 30 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M45 76 39 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M46 161 22 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M47 5 76 112 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M48 13 39 5 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M49 62 39 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29780 $Y=20590 $dt=1
M50 35 13 62 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30190 $Y=20590 $dt=1
M51 35 13 112 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M52 113 14 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M53 63 14 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=20590 $dt=1
M54 35 40 63 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=20590 $dt=1
M55 6 40 14 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M56 78 6 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M57 113 77 6 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M58 51 78 114 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M59 35 40 77 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M60 31 6 51 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M61 35 31 114 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M62 79 7 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M63 116 15 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M64 64 15 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=20590 $dt=1
M65 35 41 64 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=20590 $dt=1
M66 52 79 115 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M67 7 41 15 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M68 32 7 52 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M69 116 80 7 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M70 35 32 115 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M71 35 41 80 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M72 81 8 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M73 118 16 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M74 65 16 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=20590 $dt=1
M75 53 81 117 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M76 35 42 65 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=20590 $dt=1
M77 8 42 16 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M78 33 8 53 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=48010 $Y=800 $dt=1
M79 118 82 8 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M80 35 33 117 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=48940 $Y=800 $dt=1
M81 35 42 82 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M82 119 54 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=50070 $Y=800 $dt=1
M83 55 9 54 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=51000 $Y=800 $dt=1
M84 119 83 55 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=51930 $Y=800 $dt=1
M85 35 9 83 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=52860 $Y=800 $dt=1
M86 84 43 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M87 9 84 120 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M88 17 43 9 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M89 66 43 35 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=20590 $dt=1
M90 35 17 66 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=20590 $dt=1
M91 35 17 120 35 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
.ends WallaceFinalAdder
