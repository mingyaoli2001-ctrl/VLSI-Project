* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : FAdder                                       *
* Netlisted  : Fri Dec  5 11:51:49 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764953504730                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764953504730 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764953504730

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764953504731                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764953504731 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764953504731

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764953504732                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764953504732 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764953504732

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_764953504733                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_764953504733 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_764953504733

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_764953504735                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_764953504735 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_764953504735

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764953504730                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764953504730 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764953504730

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764953504732                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764953504732 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_764953504732

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764953504733                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764953504733 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_764953504733

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764953504734                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764953504734 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764953504734

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764953504735                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764953504735 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_764953504735

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764953504736                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764953504736 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764953504736

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764953504737                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764953504737 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=101.54 scb=0.0428868 scc=0.0113759 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764953504737

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764953504738                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764953504738 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764953504738

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764953504739                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764953504739 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764953504739

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7649535047310                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7649535047310 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7649535047310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAdder 2 6 3 9 7 8 10
** N=10 EP=7 FDC=18
X0 1 M1_PO_CDNS_764953504730 $T=1550 6040 0 90 $X=1430 $Y=5940
X1 2 M1_PO_CDNS_764953504730 $T=3090 2650 0 90 $X=2970 $Y=2550
X2 2 M1_PO_CDNS_764953504730 $T=3090 3820 0 90 $X=2970 $Y=3720
X3 2 M1_PO_CDNS_764953504730 $T=3090 4360 0 90 $X=2970 $Y=4260
X4 3 M1_PO_CDNS_764953504730 $T=3145 6870 0 90 $X=3025 $Y=6770
X5 4 M1_PO_CDNS_764953504730 $T=3720 5020 0 90 $X=3600 $Y=4920
X6 5 M2_M1_CDNS_764953504731 $T=2700 5110 0 90 $X=2570 $Y=5030
X7 4 M2_M1_CDNS_764953504731 $T=3060 2950 0 90 $X=2930 $Y=2870
X8 4 M2_M1_CDNS_764953504731 $T=3060 5520 0 90 $X=2930 $Y=5440
X9 2 M2_M1_CDNS_764953504731 $T=3450 7370 0 90 $X=3320 $Y=7290
X10 6 M2_M1_CDNS_764953504731 $T=3450 8190 0 90 $X=3320 $Y=8110
X11 2 M2_M1_CDNS_764953504731 $T=3460 3880 0 90 $X=3330 $Y=3800
X12 6 M2_M1_CDNS_764953504731 $T=4250 4700 0 90 $X=4120 $Y=4620
X13 1 M2_M1_CDNS_764953504731 $T=4700 5110 0 90 $X=4570 $Y=5030
X14 1 M2_M1_CDNS_764953504731 $T=4740 5820 0 90 $X=4610 $Y=5740
X15 5 M2_M1_CDNS_764953504731 $T=5140 5990 0 90 $X=5010 $Y=5910
X16 5 M2_M1_CDNS_764953504732 $T=2700 7470 0 90 $X=2450 $Y=7390
X17 3 M2_M1_CDNS_764953504732 $T=3820 6180 0 90 $X=3570 $Y=6100
X18 6 M2_M1_CDNS_764953504732 $T=4200 5220 0 90 $X=3950 $Y=5140
X19 6 M2_M1_CDNS_764953504732 $T=4250 4170 0 90 $X=4000 $Y=4090
X20 1 M2_M1_CDNS_764953504732 $T=4650 8090 0 90 $X=4400 $Y=8010
X21 5 M1_PO_CDNS_764953504733 $T=2700 7470 0 90 $X=2450 $Y=7370
X22 3 M1_PO_CDNS_764953504733 $T=3820 6180 0 90 $X=3570 $Y=6080
X23 6 M1_PO_CDNS_764953504733 $T=4200 5220 0 90 $X=3950 $Y=5120
X24 6 M1_PO_CDNS_764953504733 $T=4250 4170 0 90 $X=4000 $Y=4070
X25 1 M1_PO_CDNS_764953504733 $T=4650 8090 0 90 $X=4400 $Y=7990
X26 5 M1_PO_CDNS_764953504733 $T=5020 6720 0 90 $X=4770 $Y=6620
X27 3 M2_M1_CDNS_764953504735 $T=3820 2110 0 90 $X=3740 $Y=1860
X28 6 M2_M1_CDNS_764953504735 $T=4260 2110 0 90 $X=4180 $Y=1860
X29 7 4 2 nmos1v_CDNS_764953504730 $T=2220 3200 1 270 $X=1420 $Y=2690
X30 4 6 5 7 nmos1v_CDNS_764953504732 $T=2220 5270 0 90 $X=1780 $Y=5030
X31 1 3 8 7 nmos1v_CDNS_764953504732 $T=2220 6290 1 270 $X=1780 $Y=5780
X32 6 1 9 7 nmos1v_CDNS_764953504732 $T=2220 7950 0 90 $X=1780 $Y=7710
X33 1 2 6 7 nmos1v_CDNS_764953504733 $T=2220 4130 1 270 $X=1780 $Y=3620
X34 8 3 1 7 nmos1v_CDNS_764953504733 $T=2220 6610 0 90 $X=1780 $Y=6250
X35 9 3 5 7 nmos1v_CDNS_764953504733 $T=2220 7630 1 270 $X=1780 $Y=7120
X36 2 6 5 7 10 pmos1v_CDNS_764953504734 $T=5670 4040 0 90 $X=5230 $Y=3620
X37 4 6 1 7 10 pmos1v_CDNS_764953504734 $T=5670 5360 1 270 $X=5230 $Y=5030
X38 2 5 9 7 10 pmos1v_CDNS_764953504734 $T=5670 7540 0 90 $X=5230 $Y=7120
X39 3 5 8 7 10 pmos1v_CDNS_764953504735 $T=5670 6700 1 270 $X=5230 $Y=6250
X40 3 1 9 7 10 pmos1v_CDNS_764953504735 $T=5670 8040 1 270 $X=5230 $Y=7590
X41 5 6 4 7 nmos1v_CDNS_764953504736 $T=2220 4950 1 270 $X=1780 $Y=4500
X42 5 2 6 7 10 pmos1v_CDNS_764953504737 $T=5670 4540 1 270 $X=5230 $Y=4090
X43 6 1 4 7 10 pmos1v_CDNS_764953504738 $T=5670 4860 0 90 $X=5230 $Y=4500
X44 10 4 2 7 pmos1v_CDNS_764953504739 $T=5670 3200 1 270 $X=5230 $Y=2690
X45 5 3 8 7 10 pmos1v_CDNS_7649535047310 $T=5670 6200 0 90 $X=5230 $Y=5780
M0 1 6 2 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=4040 $dt=0
M1 6 2 1 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=4450 $dt=0
M2 4 6 5 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=5270 $dt=0
M3 8 3 1 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=6200 $dt=0
M4 3 1 8 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=6610 $dt=0
M5 9 5 3 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=7540 $dt=0
M6 6 1 9 7 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=7950 $dt=0
M7 5 6 2 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=5430 $Y=4040 $dt=1
M8 4 6 1 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=5430 $Y=5270 $dt=1
M9 3 5 8 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=101.512 scb=0.0428767 scc=0.0113759 $X=5430 $Y=6610 $dt=1
M10 9 5 2 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=105.522 scb=0.0482999 scc=0.011447 $X=5430 $Y=7540 $dt=1
M11 3 1 9 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=118.958 scb=0.0655284 scc=0.0136418 $X=5430 $Y=7950 $dt=1
.ends FAdder
