* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : XOR                                          *
* Netlisted  : Sun Dec  7 11:13:11 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765123987260                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765123987260 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765123987260

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765123987262                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765123987262 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765123987262

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765123987263                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765123987263 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765123987263

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765123987260                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765123987260 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765123987260

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765123987261                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765123987261 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765123987261

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR 1 2 6 5 4
** N=7 EP=5 FDC=8
X0 1 M1_PO_CDNS_765123987260 $T=320 1490 0 0 $X=220 $Y=1240
X1 2 M1_PO_CDNS_765123987260 $T=1540 2050 0 0 $X=1440 $Y=1800
X2 2 M1_PO_CDNS_765123987260 $T=3400 2050 0 0 $X=3300 $Y=1800
X3 1 M2_M1_CDNS_765123987262 $T=320 1490 0 0 $X=240 $Y=1240
X4 2 M2_M1_CDNS_765123987262 $T=1540 2050 0 0 $X=1460 $Y=1800
X5 2 M2_M1_CDNS_765123987262 $T=3400 2050 0 0 $X=3320 $Y=1800
X6 3 M2_M1_CDNS_765123987263 $T=690 3330 0 0 $X=610 $Y=3200
X7 1 M2_M1_CDNS_765123987263 $T=1190 1490 0 0 $X=1110 $Y=1360
X8 1 M2_M1_CDNS_765123987263 $T=2520 1490 0 0 $X=2440 $Y=1360
X9 3 M2_M1_CDNS_765123987263 $T=2550 3330 0 0 $X=2470 $Y=3200
X10 4 3 4 1 5 pmos1v_CDNS_765123987260 $T=420 3660 0 0 $X=0 $Y=3460
X11 1 6 4 2 5 pmos1v_CDNS_765123987260 $T=1350 3660 0 0 $X=930 $Y=3460
X12 3 6 4 7 5 pmos1v_CDNS_765123987260 $T=2370 3660 1 180 $X=1860 $Y=3460
X13 4 7 4 2 5 pmos1v_CDNS_765123987260 $T=3300 3660 1 180 $X=2790 $Y=3460
X14 5 5 1 3 nmos1v_CDNS_765123987261 $T=420 800 0 0 $X=0 $Y=240
X15 6 5 2 3 nmos1v_CDNS_765123987261 $T=1440 800 1 180 $X=930 $Y=240
X16 6 5 7 1 nmos1v_CDNS_765123987261 $T=2280 800 0 0 $X=1860 $Y=240
X17 5 5 2 7 nmos1v_CDNS_765123987261 $T=3300 800 1 180 $X=2790 $Y=240
M0 3 1 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=420 $Y=3660 $dt=1
M1 6 2 1 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1350 $Y=3660 $dt=1
M2 3 7 6 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2280 $Y=3660 $dt=1
M3 4 2 7 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3210 $Y=3660 $dt=1
.ends XOR
