* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : XORgate                                      *
* Netlisted  : Mon Oct 20 22:25:27 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_761013523105                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_761013523105 1 2 3 5
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=4.5e-07 sca=112.466 scb=0.0581753 scc=0.0119018 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_761013523105

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523106                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523106 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.55e-07 sca=6.629 scb=0.00319937 scc=2.08619e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_761013523106

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523107                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523107 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=4.5e-07 sb=2.45e-07 sca=7.61443 scb=0.00488365 scc=5.56751e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_761013523107

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523108                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523108 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.55e-07 sca=7.61443 scb=0.00488365 scc=5.56751e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_761013523108

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XORgate                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XORgate a b gnd vdd y
** N=11 EP=5 FDC=12
X21 y 6 8 vdd pmos1v_CDNS_761013523105 $T=5440 -2790 1 180 $X=4990 $Y=-2990
X22 gnd 6 10 nmos1v_CDNS_761013523106 $T=5650 -4060 1 180 $X=5360 $Y=-4260
X23 y a 11 gnd nmos1v_CDNS_761013523107 $T=5030 -4060 1 180 $X=4740 $Y=-4260
X24 gnd b 11 nmos1v_CDNS_761013523108 $T=4730 -4060 0 0 $X=4310 $Y=-4260
M0 6 b gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=5.97505 scb=0.00216741 scc=8.45511e-06 $X=1110 $Y=-4080 $dt=0
M1 5 a gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.629 scb=0.00319937 scc=2.08619e-05 $X=3020 $Y=-4070 $dt=0
M2 10 5 y gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=4.5e-07 sb=2.45e-07 sca=6.629 scb=0.00319937 scc=2.08619e-05 $X=5350 $Y=-4060 $dt=0
M3 6 b vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=133.279 scb=0.0807128 scc=0.0160465 $X=1110 $Y=-2710 $dt=1
M4 5 a vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=132.037 scb=0.0810715 scc=0.0154938 $X=3020 $Y=-2800 $dt=1
M5 7 5 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.55e-07 sca=65.2428 scb=0.0627023 scc=0.00830595 $X=4730 $Y=-2790 $dt=1
M6 y b 7 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=4.5e-07 sca=56.4563 scb=0.0530432 scc=0.0064557 $X=4940 $Y=-2790 $dt=1
M7 vdd a 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=5.55e-07 sb=1.4e-07 sca=119.893 scb=0.0639272 scc=0.0138773 $X=5560 $Y=-2790 $dt=1
.ends XORgate
