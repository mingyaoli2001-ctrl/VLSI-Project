* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : XORgate                                      *
* Netlisted  : Mon Oct 20 22:25:27 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_NWELL_CDNS_761013523100                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_NWELL_CDNS_761013523100 1
** N=1 EP=1 FDC=0
.ends M1_NWELL_CDNS_761013523100

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PSUB_CDNS_761013523101                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PSUB_CDNS_761013523101 1
** N=1 EP=1 FDC=0
.ends M1_PSUB_CDNS_761013523101

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_761013523102                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_761013523102 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_761013523102

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_761013523103                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_761013523103 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_761013523103

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_761013523100                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_761013523100 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_761013523100

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523101                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523101 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_761013523101

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_761013523104                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_761013523104 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_761013523104

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_761013523105                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_761013523105 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=4.5e-07 sca=112.466 scb=0.0581753 scc=0.0119018 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_761013523105

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523106                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523106 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.55e-07 sca=6.629 scb=0.00319937 scc=2.08619e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_761013523106

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523107                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523107 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=4.5e-07 sb=2.45e-07 sca=7.61443 scb=0.00488365 scc=5.56751e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_761013523107

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_761013523108                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_761013523108 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.55e-07 sca=7.61443 scb=0.00488365 scc=5.56751e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_761013523108

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XORgate                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XORgate 4 3 2 1 9
** N=11 EP=5 FDC=12
X0 1 M1_NWELL_CDNS_761013523100 $T=950 -1770 0 0 $X=630 $Y=-2090
X1 1 M1_NWELL_CDNS_761013523100 $T=2860 -1880 0 0 $X=2540 $Y=-2200
X2 1 M1_NWELL_CDNS_761013523100 $T=5810 -2040 0 0 $X=5490 $Y=-2360
X3 2 M1_PSUB_CDNS_761013523101 $T=950 -4880 0 0 $X=730 $Y=-5100
X4 2 M1_PSUB_CDNS_761013523101 $T=2860 -4880 0 0 $X=2640 $Y=-5100
X5 2 M1_PSUB_CDNS_761013523101 $T=4570 -5240 0 0 $X=4350 $Y=-5460
X6 3 M1_PO_CDNS_761013523102 $T=560 -3270 0 0 $X=460 $Y=-3390
X7 4 M1_PO_CDNS_761013523102 $T=2500 -3270 0 0 $X=2400 $Y=-3390
X8 5 M1_PO_CDNS_761013523102 $T=3760 -2020 0 0 $X=3660 $Y=-2140
X9 6 M1_PO_CDNS_761013523102 $T=5260 -1700 0 0 $X=5160 $Y=-1820
X10 5 M1_PO_CDNS_761013523102 $T=5410 -4830 0 0 $X=5310 $Y=-4950
X11 6 M2_M1_CDNS_761013523103 $T=1370 -1060 0 0 $X=1290 $Y=-1190
X12 5 M2_M1_CDNS_761013523103 $T=3700 -4830 0 0 $X=3620 $Y=-4960
X13 5 M2_M1_CDNS_761013523103 $T=4950 -4830 0 0 $X=4870 $Y=-4960
X14 6 M2_M1_CDNS_761013523103 $T=5260 -1060 0 0 $X=5180 $Y=-1190
X15 1 6 3 2 pmos1v_CDNS_761013523100 $T=1110 -2710 0 0 $X=690 $Y=-2910
X16 1 5 4 2 pmos1v_CDNS_761013523100 $T=3020 -2800 0 0 $X=2600 $Y=-3000
X17 2 6 3 nmos1v_CDNS_761013523101 $T=1110 -4080 0 0 $X=690 $Y=-4280
X18 2 5 4 nmos1v_CDNS_761013523101 $T=3020 -4070 0 0 $X=2600 $Y=-4270
X19 1 5 7 2 pmos1v_CDNS_761013523104 $T=4730 -2790 0 0 $X=4310 $Y=-2990
X20 1 4 8 2 pmos1v_CDNS_761013523104 $T=5650 -2550 0 180 $X=5360 $Y=-2990
X21 9 6 8 2 1 pmos1v_CDNS_761013523105 $T=5440 -2790 1 180 $X=4990 $Y=-2990
X22 2 6 10 nmos1v_CDNS_761013523106 $T=5650 -4060 1 180 $X=5360 $Y=-4260
X23 9 4 11 2 nmos1v_CDNS_761013523107 $T=5030 -4060 1 180 $X=4740 $Y=-4260
X24 2 3 11 nmos1v_CDNS_761013523108 $T=4730 -4060 0 0 $X=4310 $Y=-4260
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=5.97505 scb=0.00216741 scc=8.45511e-06 $X=1110 $Y=-4080 $dt=0
M1 5 4 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.629 scb=0.00319937 scc=2.08619e-05 $X=3020 $Y=-4070 $dt=0
M2 10 5 9 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=4.5e-07 sb=2.45e-07 sca=6.629 scb=0.00319937 scc=2.08619e-05 $X=5350 $Y=-4060 $dt=0
M3 6 3 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=133.279 scb=0.0807128 scc=0.0160465 $X=1110 $Y=-2710 $dt=1
M4 5 4 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=132.037 scb=0.0810715 scc=0.0154938 $X=3020 $Y=-2800 $dt=1
M5 7 5 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=5.55e-07 sca=65.2428 scb=0.0627023 scc=0.00830595 $X=4730 $Y=-2790 $dt=1
M6 9 3 7 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=4.5e-07 sca=56.4563 scb=0.0530432 scc=0.0064557 $X=4940 $Y=-2790 $dt=1
M7 1 4 8 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=5.55e-07 sb=1.4e-07 sca=119.893 scb=0.0639272 scc=0.0138773 $X=5560 $Y=-2790 $dt=1
.ends XORgate
