* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : WallaceMultiplier                            *
* Netlisted  : Thu Dec  4 17:53:32 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceMultiplier                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceMultiplier a<0> a<1> a<2> a<3> a<4> a<5> a<6> a<7> b<0> b<1>
+ b<2> b<3> b<4> b<5> b<6> b<7> gnd p00 p01 p02
+ p03 p04 p05 p06 p07 p10 p11 p12 p13 p14
+ p15 p16 p17 p20 p21 p22 p23 p24 p25 p26
+ p27 p30 p31 p32 p33 p34 p35 p36 p37 p40
+ p41 p42 p43 p44 p45 p46 p47 p50 p51 p52
+ p53 p54 p55 p56 p57 p60 p61 p62 p63 p64
+ p65 p66 p67 p70 p71 p72 p73 p74 p75 p76
+ p77 vdd
** N=210 EP=82 FDC=384
M0 147 a<7> 83 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=33350 $dt=0
M1 148 a<6> 84 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=34150 $dt=0
M2 149 a<5> 85 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=37890 $dt=0
M3 150 a<4> 86 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=38690 $dt=0
M4 151 a<3> 87 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=42430 $dt=0
M5 152 a<2> 88 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=43230 $dt=0
M6 153 a<1> 89 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=46970 $dt=0
M7 154 a<0> 90 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=47770 $dt=0
M8 gnd b<0> 147 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=33350 $dt=0
M9 gnd b<0> 148 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=34150 $dt=0
M10 gnd b<0> 149 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=37890 $dt=0
M11 gnd b<0> 150 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=38690 $dt=0
M12 gnd b<0> 151 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=42430 $dt=0
M13 gnd b<0> 152 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=43230 $dt=0
M14 gnd b<0> 153 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=46970 $dt=0
M15 gnd b<0> 154 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=47770 $dt=0
M16 p07 83 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=33360 $dt=0
M17 p06 84 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=34140 $dt=0
M18 p05 85 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=37900 $dt=0
M19 p04 86 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=38680 $dt=0
M20 p03 87 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=42440 $dt=0
M21 p02 88 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=43220 $dt=0
M22 p01 89 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=46980 $dt=0
M23 p00 90 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=47760 $dt=0
M24 155 a<7> 91 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=33340 $dt=0
M25 156 a<6> 92 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=34140 $dt=0
M26 157 a<5> 93 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=37890 $dt=0
M27 158 a<4> 94 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=38690 $dt=0
M28 159 a<3> 95 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=42430 $dt=0
M29 160 a<2> 96 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=43230 $dt=0
M30 161 a<1> 97 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=46970 $dt=0
M31 162 a<0> 98 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=47770 $dt=0
M32 gnd b<1> 155 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=33340 $dt=0
M33 gnd b<1> 156 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=34140 $dt=0
M34 gnd b<1> 157 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=37890 $dt=0
M35 gnd b<1> 158 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=38690 $dt=0
M36 gnd b<1> 159 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=42430 $dt=0
M37 gnd b<1> 160 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=43230 $dt=0
M38 gnd b<1> 161 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=46970 $dt=0
M39 gnd b<1> 162 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=47770 $dt=0
M40 p17 91 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=33350 $dt=0
M41 p16 92 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=34130 $dt=0
M42 p15 93 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=37900 $dt=0
M43 p14 94 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=38680 $dt=0
M44 p13 95 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=42440 $dt=0
M45 p12 96 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=43220 $dt=0
M46 p11 97 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=46980 $dt=0
M47 p10 98 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=47760 $dt=0
M48 163 a<7> 99 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=33340 $dt=0
M49 164 a<6> 100 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=34140 $dt=0
M50 165 a<5> 101 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=37890 $dt=0
M51 166 a<4> 102 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=38690 $dt=0
M52 167 a<3> 103 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=42430 $dt=0
M53 168 a<2> 104 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=43230 $dt=0
M54 169 a<1> 105 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=46970 $dt=0
M55 170 a<0> 106 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=47770 $dt=0
M56 gnd b<2> 163 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=33340 $dt=0
M57 gnd b<2> 164 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=34140 $dt=0
M58 gnd b<2> 165 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=37890 $dt=0
M59 gnd b<2> 166 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=38690 $dt=0
M60 gnd b<2> 167 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=42430 $dt=0
M61 gnd b<2> 168 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=43230 $dt=0
M62 gnd b<2> 169 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=46970 $dt=0
M63 gnd b<2> 170 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=47770 $dt=0
M64 p27 99 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=33350 $dt=0
M65 p26 100 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=34130 $dt=0
M66 p25 101 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=37900 $dt=0
M67 p24 102 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=38680 $dt=0
M68 p23 103 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=42440 $dt=0
M69 p22 104 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=43220 $dt=0
M70 p21 105 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=46980 $dt=0
M71 p20 106 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=47760 $dt=0
M72 171 a<7> 107 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=33340 $dt=0
M73 172 a<6> 108 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=34140 $dt=0
M74 173 a<5> 109 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=37890 $dt=0
M75 174 a<4> 110 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=38690 $dt=0
M76 175 a<3> 111 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=42430 $dt=0
M77 176 a<2> 112 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=43230 $dt=0
M78 177 a<1> 113 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=46970 $dt=0
M79 178 a<0> 114 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=47770 $dt=0
M80 gnd b<3> 171 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=33340 $dt=0
M81 gnd b<3> 172 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=34140 $dt=0
M82 gnd b<3> 173 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=37890 $dt=0
M83 gnd b<3> 174 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=38690 $dt=0
M84 gnd b<3> 175 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=42430 $dt=0
M85 gnd b<3> 176 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=43230 $dt=0
M86 gnd b<3> 177 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=46970 $dt=0
M87 gnd b<3> 178 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=47770 $dt=0
M88 p37 107 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=33350 $dt=0
M89 p36 108 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=34130 $dt=0
M90 p35 109 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=37900 $dt=0
M91 p34 110 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=38680 $dt=0
M92 p33 111 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=42440 $dt=0
M93 p32 112 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=43220 $dt=0
M94 p31 113 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=46980 $dt=0
M95 p30 114 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=47760 $dt=0
M96 179 a<7> 115 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=33340 $dt=0
M97 180 a<6> 116 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=34140 $dt=0
M98 181 a<5> 117 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=37890 $dt=0
M99 182 a<4> 118 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=38690 $dt=0
M100 183 a<3> 119 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=42430 $dt=0
M101 184 a<2> 120 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=43230 $dt=0
M102 185 a<1> 121 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=46970 $dt=0
M103 186 a<0> 122 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=47770 $dt=0
M104 gnd b<4> 179 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=33340 $dt=0
M105 gnd b<4> 180 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=34140 $dt=0
M106 gnd b<4> 181 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=37890 $dt=0
M107 gnd b<4> 182 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=38690 $dt=0
M108 gnd b<4> 183 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=42430 $dt=0
M109 gnd b<4> 184 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=43230 $dt=0
M110 gnd b<4> 185 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=46970 $dt=0
M111 gnd b<4> 186 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=47770 $dt=0
M112 p47 115 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=33350 $dt=0
M113 p46 116 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=34130 $dt=0
M114 p45 117 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=37900 $dt=0
M115 p44 118 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=38680 $dt=0
M116 p43 119 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=42440 $dt=0
M117 p42 120 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=43220 $dt=0
M118 p41 121 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=46980 $dt=0
M119 p40 122 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=47760 $dt=0
M120 187 a<7> 123 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=33340 $dt=0
M121 188 a<6> 124 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=34140 $dt=0
M122 189 a<5> 125 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=37890 $dt=0
M123 190 a<4> 126 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=38690 $dt=0
M124 191 a<3> 127 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=42430 $dt=0
M125 192 a<2> 128 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=43230 $dt=0
M126 193 a<1> 129 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=46970 $dt=0
M127 194 a<0> 130 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=47770 $dt=0
M128 gnd b<5> 187 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=33340 $dt=0
M129 gnd b<5> 188 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=34140 $dt=0
M130 gnd b<5> 189 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=37890 $dt=0
M131 gnd b<5> 190 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=38690 $dt=0
M132 gnd b<5> 191 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=42430 $dt=0
M133 gnd b<5> 192 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=43230 $dt=0
M134 gnd b<5> 193 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=46970 $dt=0
M135 gnd b<5> 194 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=47770 $dt=0
M136 p57 123 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=33350 $dt=0
M137 p56 124 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=34130 $dt=0
M138 p55 125 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=37900 $dt=0
M139 p54 126 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=38680 $dt=0
M140 p53 127 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=42440 $dt=0
M141 p52 128 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=43220 $dt=0
M142 p51 129 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=46980 $dt=0
M143 p50 130 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=47760 $dt=0
M144 195 a<7> 131 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=33350 $dt=0
M145 196 a<6> 132 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=34140 $dt=0
M146 197 a<5> 133 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=37890 $dt=0
M147 198 a<4> 134 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=38690 $dt=0
M148 199 a<3> 135 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=42430 $dt=0
M149 200 a<2> 136 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=43230 $dt=0
M150 201 a<1> 137 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=46970 $dt=0
M151 202 a<0> 138 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=47770 $dt=0
M152 gnd b<6> 195 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=33350 $dt=0
M153 gnd b<6> 196 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=34140 $dt=0
M154 gnd b<6> 197 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=37890 $dt=0
M155 gnd b<6> 198 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=38690 $dt=0
M156 gnd b<6> 199 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=42430 $dt=0
M157 gnd b<6> 200 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=43230 $dt=0
M158 gnd b<6> 201 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=46970 $dt=0
M159 gnd b<6> 202 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=47770 $dt=0
M160 p67 131 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=33360 $dt=0
M161 p66 132 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=34130 $dt=0
M162 p65 133 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=37900 $dt=0
M163 p64 134 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=38680 $dt=0
M164 p63 135 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=42440 $dt=0
M165 p62 136 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=43220 $dt=0
M166 p61 137 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=46980 $dt=0
M167 p60 138 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=47760 $dt=0
M168 203 a<7> 139 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=33350 $dt=0
M169 204 a<6> 140 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=34150 $dt=0
M170 205 a<5> 141 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=37890 $dt=0
M171 206 a<4> 142 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=38690 $dt=0
M172 207 a<3> 143 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=42430 $dt=0
M173 208 a<2> 144 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=43230 $dt=0
M174 209 a<1> 145 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=46970 $dt=0
M175 210 a<0> 146 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=47770 $dt=0
M176 gnd b<7> 203 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=33350 $dt=0
M177 gnd b<7> 204 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=34150 $dt=0
M178 gnd b<7> 205 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=37890 $dt=0
M179 gnd b<7> 206 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=38690 $dt=0
M180 gnd b<7> 207 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=42430 $dt=0
M181 gnd b<7> 208 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=43230 $dt=0
M182 gnd b<7> 209 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=46970 $dt=0
M183 gnd b<7> 210 gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=47770 $dt=0
M184 p77 139 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=33360 $dt=0
M185 p76 140 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=34140 $dt=0
M186 p75 141 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=37900 $dt=0
M187 p74 142 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=38680 $dt=0
M188 p73 143 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=42440 $dt=0
M189 p72 144 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=43220 $dt=0
M190 p71 145 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=46980 $dt=0
M191 p70 146 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=47760 $dt=0
M192 83 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=31910 $dt=1
M193 84 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=35590 $dt=1
M194 85 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=36450 $dt=1
M195 86 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40130 $dt=1
M196 87 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40990 $dt=1
M197 88 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=44670 $dt=1
M198 89 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=45530 $dt=1
M199 90 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=49210 $dt=1
M200 vdd b<0> 83 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=31910 $dt=1
M201 vdd b<0> 84 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=35590 $dt=1
M202 vdd b<0> 85 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=36450 $dt=1
M203 vdd b<0> 86 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40130 $dt=1
M204 vdd b<0> 87 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40990 $dt=1
M205 vdd b<0> 88 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=44670 $dt=1
M206 vdd b<0> 89 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=45530 $dt=1
M207 vdd b<0> 90 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=49210 $dt=1
M208 p07 83 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=31860 $dt=1
M209 p06 84 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=35400 $dt=1
M210 p05 85 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=36400 $dt=1
M211 p04 86 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=39940 $dt=1
M212 p03 87 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=40940 $dt=1
M213 p02 88 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=44480 $dt=1
M214 p01 89 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=45480 $dt=1
M215 p00 90 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=49020 $dt=1
M216 91 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=31900 $dt=1
M217 92 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=35580 $dt=1
M218 93 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=36450 $dt=1
M219 94 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40130 $dt=1
M220 95 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40990 $dt=1
M221 96 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=44670 $dt=1
M222 97 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=45530 $dt=1
M223 98 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=49210 $dt=1
M224 vdd b<1> 91 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=31900 $dt=1
M225 vdd b<1> 92 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=35580 $dt=1
M226 vdd b<1> 93 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=36450 $dt=1
M227 vdd b<1> 94 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40130 $dt=1
M228 vdd b<1> 95 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40990 $dt=1
M229 vdd b<1> 96 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=44670 $dt=1
M230 vdd b<1> 97 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=45530 $dt=1
M231 vdd b<1> 98 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=49210 $dt=1
M232 p17 91 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=31850 $dt=1
M233 p16 92 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=35390 $dt=1
M234 p15 93 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=36400 $dt=1
M235 p14 94 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=39940 $dt=1
M236 p13 95 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=40940 $dt=1
M237 p12 96 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=44480 $dt=1
M238 p11 97 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=45480 $dt=1
M239 p10 98 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=49020 $dt=1
M240 99 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=31900 $dt=1
M241 100 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=35580 $dt=1
M242 101 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=36450 $dt=1
M243 102 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40130 $dt=1
M244 103 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40990 $dt=1
M245 104 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=44670 $dt=1
M246 105 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=45530 $dt=1
M247 106 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=49210 $dt=1
M248 vdd b<2> 99 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=31900 $dt=1
M249 vdd b<2> 100 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=35580 $dt=1
M250 vdd b<2> 101 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=36450 $dt=1
M251 vdd b<2> 102 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40130 $dt=1
M252 vdd b<2> 103 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40990 $dt=1
M253 vdd b<2> 104 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=44670 $dt=1
M254 vdd b<2> 105 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=45530 $dt=1
M255 vdd b<2> 106 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=49210 $dt=1
M256 p27 99 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=31850 $dt=1
M257 p26 100 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=35390 $dt=1
M258 p25 101 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=36400 $dt=1
M259 p24 102 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=39940 $dt=1
M260 p23 103 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=40940 $dt=1
M261 p22 104 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=44480 $dt=1
M262 p21 105 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=45480 $dt=1
M263 p20 106 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=49020 $dt=1
M264 107 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=31900 $dt=1
M265 108 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=35580 $dt=1
M266 109 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=36450 $dt=1
M267 110 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40130 $dt=1
M268 111 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40990 $dt=1
M269 112 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=44670 $dt=1
M270 113 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=45530 $dt=1
M271 114 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=49210 $dt=1
M272 vdd b<3> 107 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=31900 $dt=1
M273 vdd b<3> 108 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=35580 $dt=1
M274 vdd b<3> 109 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=36450 $dt=1
M275 vdd b<3> 110 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40130 $dt=1
M276 vdd b<3> 111 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40990 $dt=1
M277 vdd b<3> 112 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=44670 $dt=1
M278 vdd b<3> 113 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=45530 $dt=1
M279 vdd b<3> 114 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=49210 $dt=1
M280 p37 107 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=31850 $dt=1
M281 p36 108 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=35390 $dt=1
M282 p35 109 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=36400 $dt=1
M283 p34 110 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=39940 $dt=1
M284 p33 111 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=40940 $dt=1
M285 p32 112 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=44480 $dt=1
M286 p31 113 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=45480 $dt=1
M287 p30 114 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=49020 $dt=1
M288 115 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=31900 $dt=1
M289 116 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=35580 $dt=1
M290 117 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=36450 $dt=1
M291 118 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40130 $dt=1
M292 119 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40990 $dt=1
M293 120 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=44670 $dt=1
M294 121 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=45530 $dt=1
M295 122 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=49210 $dt=1
M296 vdd b<4> 115 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=31900 $dt=1
M297 vdd b<4> 116 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=35580 $dt=1
M298 vdd b<4> 117 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=36450 $dt=1
M299 vdd b<4> 118 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40130 $dt=1
M300 vdd b<4> 119 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40990 $dt=1
M301 vdd b<4> 120 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=44670 $dt=1
M302 vdd b<4> 121 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=45530 $dt=1
M303 vdd b<4> 122 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=49210 $dt=1
M304 p47 115 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=31850 $dt=1
M305 p46 116 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=35390 $dt=1
M306 p45 117 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=36400 $dt=1
M307 p44 118 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=39940 $dt=1
M308 p43 119 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=40940 $dt=1
M309 p42 120 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=44480 $dt=1
M310 p41 121 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=45480 $dt=1
M311 p40 122 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=49020 $dt=1
M312 123 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=31900 $dt=1
M313 124 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=35580 $dt=1
M314 125 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=36450 $dt=1
M315 126 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40130 $dt=1
M316 127 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40990 $dt=1
M317 128 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=44670 $dt=1
M318 129 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=45530 $dt=1
M319 130 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=49210 $dt=1
M320 vdd b<5> 123 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=31900 $dt=1
M321 vdd b<5> 124 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=35580 $dt=1
M322 vdd b<5> 125 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=36450 $dt=1
M323 vdd b<5> 126 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40130 $dt=1
M324 vdd b<5> 127 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40990 $dt=1
M325 vdd b<5> 128 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=44670 $dt=1
M326 vdd b<5> 129 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=45530 $dt=1
M327 vdd b<5> 130 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=49210 $dt=1
M328 p57 123 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=31850 $dt=1
M329 p56 124 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=35390 $dt=1
M330 p55 125 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=36400 $dt=1
M331 p54 126 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=39940 $dt=1
M332 p53 127 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=40940 $dt=1
M333 p52 128 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=44480 $dt=1
M334 p51 129 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=45480 $dt=1
M335 p50 130 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=49020 $dt=1
M336 131 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=31910 $dt=1
M337 132 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=35580 $dt=1
M338 133 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=36450 $dt=1
M339 134 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40130 $dt=1
M340 135 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40990 $dt=1
M341 136 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=44670 $dt=1
M342 137 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=45530 $dt=1
M343 138 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=49210 $dt=1
M344 vdd b<6> 131 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=31910 $dt=1
M345 vdd b<6> 132 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=35580 $dt=1
M346 vdd b<6> 133 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=36450 $dt=1
M347 vdd b<6> 134 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40130 $dt=1
M348 vdd b<6> 135 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40990 $dt=1
M349 vdd b<6> 136 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=44670 $dt=1
M350 vdd b<6> 137 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=45530 $dt=1
M351 vdd b<6> 138 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=49210 $dt=1
M352 p67 131 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=31860 $dt=1
M353 p66 132 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=35390 $dt=1
M354 p65 133 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=36400 $dt=1
M355 p64 134 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=39940 $dt=1
M356 p63 135 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=40940 $dt=1
M357 p62 136 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=44480 $dt=1
M358 p61 137 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=45480 $dt=1
M359 p60 138 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=49020 $dt=1
M360 139 a<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=31910 $dt=1
M361 140 a<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=35590 $dt=1
M362 141 a<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=36450 $dt=1
M363 142 a<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40130 $dt=1
M364 143 a<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40990 $dt=1
M365 144 a<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=44670 $dt=1
M366 145 a<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=45530 $dt=1
M367 146 a<0> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=49210 $dt=1
M368 vdd b<7> 139 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=31910 $dt=1
M369 vdd b<7> 140 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=35590 $dt=1
M370 vdd b<7> 141 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=36450 $dt=1
M371 vdd b<7> 142 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40130 $dt=1
M372 vdd b<7> 143 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40990 $dt=1
M373 vdd b<7> 144 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=44670 $dt=1
M374 vdd b<7> 145 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=45530 $dt=1
M375 vdd b<7> 146 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=49210 $dt=1
M376 p77 139 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=31860 $dt=1
M377 p76 140 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=35400 $dt=1
M378 p75 141 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=36400 $dt=1
M379 p74 142 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=39940 $dt=1
M380 p73 143 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=40940 $dt=1
M381 p72 144 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=44480 $dt=1
M382 p71 145 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=45480 $dt=1
M383 p70 146 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=49020 $dt=1
.ends WallaceMultiplier
