* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : WallaceProject                               *
* Netlisted  : Fri Dec 12 21:35:11 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765593305580                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765593305580 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765593305580

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765593305581                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765593305581 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765593305581

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765593305582                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765593305582 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765593305582

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765593305583                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765593305583 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765593305583

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765593305584                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765593305584 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765593305584

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765593305585                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765593305585 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765593305585

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765593305586                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765593305586 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765593305586

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765593305587                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765593305587 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765593305587

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765593305588                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765593305588 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765593305588

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765593305589                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765593305589 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765593305589

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055810                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055810 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055811                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055811 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055812                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055812 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055813                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055813 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055814                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055814 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055815                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055815 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055816                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055816 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055817                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055817 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055818                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055818 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055820                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055820 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055821                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055821 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055821

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055822                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055822 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055822

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055823                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055823 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055823

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055824                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055824 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055824

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055825                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055825 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055825

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055828                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055828 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055828

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055829                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055829 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055829

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055830                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055830 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055830

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055831                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055831 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055831

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055832                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055832 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055832

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055833                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055833 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055833

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055836                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055836 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055836

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055838                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055838 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055838

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7655933055841                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7655933055841 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7655933055841

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765593305580                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765593305580 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765593305580

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765593305581                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765593305581 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765593305581

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: Diver                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt Diver 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
X0 1 M1_PO_CDNS_7655933055841 $T=1260 -2440 0 0 $X=1160 $Y=-2560
X1 5 M1_PO_CDNS_7655933055841 $T=2200 -2440 0 0 $X=2100 $Y=-2560
X2 2 2 1 5 3 pmos1v_CDNS_765593305580 $T=1340 -2060 0 0 $X=920 $Y=-2260
X3 2 2 5 4 3 pmos1v_CDNS_765593305580 $T=2270 -2060 0 0 $X=1850 $Y=-2260
X4 3 3 1 5 nmos1v_CDNS_765593305581 $T=1340 -3070 0 0 $X=920 $Y=-3630
X5 3 3 5 4 nmos1v_CDNS_765593305581 $T=2270 -3070 0 0 $X=1850 $Y=-3630
.ends Diver

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055843                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055843 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055843

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7655933055844                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7655933055844 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7655933055844

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055845                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055845 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055845

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7655933055846                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7655933055846 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7655933055846

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765593305582                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765593305582 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765593305582

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765593305583                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765593305583 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765593305583

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765593305584                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765593305584 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765593305584

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765593305585                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765593305585 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765593305585

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765593305586                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765593305586 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765593305586

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765593305587                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765593305587 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765593305587

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765593305588                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765593305588 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765593305588

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765593305589                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765593305589 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765593305589

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055810                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055810 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7655933055810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055811                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055811 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7655933055811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055812                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055812 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7655933055812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=8
X0 1 M2_M1_CDNS_765593305586 $T=2220 -7390 0 90 $X=2090 $Y=-7470
X1 1 M2_M1_CDNS_765593305586 $T=2220 -4680 0 90 $X=2090 $Y=-4760
X2 7 M2_M1_CDNS_765593305586 $T=4200 -2840 0 90 $X=4070 $Y=-2920
X3 8 M2_M1_CDNS_765593305586 $T=4570 -3920 0 90 $X=4440 $Y=-4000
X4 9 M2_M1_CDNS_765593305588 $T=1300 -5710 0 90 $X=1170 $Y=-5840
X5 9 M2_M1_CDNS_765593305588 $T=1300 -4270 0 90 $X=1170 $Y=-4400
X6 6 6 4 8 2 pmos1v_CDNS_765593305580 $T=5520 -3500 0 270 $X=5320 $Y=-4010
X7 6 6 5 7 2 pmos1v_CDNS_765593305580 $T=5520 -2570 0 270 $X=5320 $Y=-3080
X8 2 2 4 8 nmos1v_CDNS_765593305581 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X9 2 2 5 7 nmos1v_CDNS_765593305581 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X10 8 M2_M1_CDNS_7655933055843 $T=2340 -4370 0 90 $X=2090 $Y=-4450
X11 8 M2_M1_CDNS_7655933055843 $T=2930 -6480 0 90 $X=2680 $Y=-6560
X12 8 M2_M1_CDNS_7655933055843 $T=2950 -5710 0 90 $X=2700 $Y=-5790
X13 4 M2_M1_CDNS_7655933055843 $T=3490 -4140 0 90 $X=3240 $Y=-4220
X14 4 M2_M1_CDNS_7655933055843 $T=3500 -3460 0 90 $X=3250 $Y=-3540
X15 10 M2_M1_CDNS_7655933055843 $T=5640 -5920 0 90 $X=5390 $Y=-6000
X16 10 M2_M1_CDNS_7655933055843 $T=5640 -5080 0 90 $X=5390 $Y=-5160
X17 10 M2_M1_CDNS_7655933055843 $T=5640 -4300 0 90 $X=5390 $Y=-4380
X18 8 M1_PO_CDNS_7655933055844 $T=2340 -4370 0 90 $X=2090 $Y=-4470
X19 8 M1_PO_CDNS_7655933055844 $T=2930 -6480 0 90 $X=2680 $Y=-6580
X20 8 M1_PO_CDNS_7655933055844 $T=2950 -5710 0 90 $X=2700 $Y=-5810
X21 4 M1_PO_CDNS_7655933055844 $T=3490 -4140 0 90 $X=3240 $Y=-4240
X22 4 M1_PO_CDNS_7655933055844 $T=3500 -3460 0 90 $X=3250 $Y=-3560
X23 4 M2_M1_CDNS_7655933055845 $T=3500 -4810 0 0 $X=3250 $Y=-4940
X24 4 M2_M1_CDNS_7655933055845 $T=3500 -1930 0 0 $X=3250 $Y=-2060
X25 7 M2_M1_CDNS_7655933055845 $T=4210 -6730 0 0 $X=3960 $Y=-6860
X26 7 M2_M1_CDNS_7655933055845 $T=4210 -5370 0 0 $X=3960 $Y=-5500
X27 8 M2_M1_CDNS_7655933055845 $T=4540 -5740 0 0 $X=4290 $Y=-5870
X28 5 M2_M1_CDNS_7655933055845 $T=4960 -4960 0 0 $X=4710 $Y=-5090
X29 5 M2_M1_CDNS_7655933055845 $T=4960 -2500 0 0 $X=4710 $Y=-2630
X30 4 M1_PO_CDNS_7655933055846 $T=3500 -4810 0 0 $X=3260 $Y=-4910
X31 7 M1_PO_CDNS_7655933055846 $T=4210 -6730 0 0 $X=3970 $Y=-6830
X32 7 M1_PO_CDNS_7655933055846 $T=4210 -5370 0 0 $X=3970 $Y=-5470
X33 8 M1_PO_CDNS_7655933055846 $T=4540 -5740 0 0 $X=4300 $Y=-5840
X34 5 M1_PO_CDNS_7655933055846 $T=4960 -4960 0 0 $X=4720 $Y=-5060
X35 5 M1_PO_CDNS_7655933055846 $T=4960 -2500 0 0 $X=4720 $Y=-2600
X36 1 5 10 2 6 pmos1v_CDNS_765593305582 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 2 7 3 nmos1v_CDNS_765593305583 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 10 6 7 2 pmos1v_CDNS_765593305584 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 6 8 11 2 pmos1v_CDNS_765593305585 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 3 7 11 2 6 pmos1v_CDNS_765593305586 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X41 2 3 8 2 nmos1v_CDNS_765593305587 $T=1570 -6390 0 270 $X=1370 $Y=-6840
X42 9 1 8 2 nmos1v_CDNS_765593305587 $T=1570 -4430 0 270 $X=1370 $Y=-4880
X43 9 7 2 2 nmos1v_CDNS_765593305588 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 4 1 12 2 nmos1v_CDNS_765593305589 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 2 5 12 nmos1v_CDNS_7655933055810 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 10 8 6 2 pmos1v_CDNS_7655933055811 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 10 4 1 2 6 pmos1v_CDNS_7655933055812 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 2 8 3 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 2 7 9 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=6.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-5550 $dt=0
M2 9 8 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M3 2 4 8 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-3590 $dt=0
M4 2 5 7 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1580 $Y=-2660 $dt=0
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055813                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055813 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_7655933055813

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055814                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055814 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7655933055814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055815                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055815 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_7655933055815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055816                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055816 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7655933055816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055817                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055817 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7655933055817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055818                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055818 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7655933055818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=0
X0 5 M3_M2_CDNS_765593305585 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X1 1 M2_M1_CDNS_765593305586 $T=1510 -2070 0 0 $X=1430 $Y=-2200
X2 1 M2_M1_CDNS_765593305586 $T=3010 -2070 0 0 $X=2930 $Y=-2200
X3 5 M2_M1_CDNS_7655933055829 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X4 2 M1_PO_CDNS_7655933055841 $T=1870 -1670 0 0 $X=1770 $Y=-1790
X5 1 M1_PO_CDNS_7655933055841 $T=2510 -2070 0 0 $X=2410 $Y=-2190
X6 6 M1_PO_CDNS_7655933055841 $T=4500 -2020 0 0 $X=4400 $Y=-2140
X7 4 5 6 nmos1v_CDNS_7655933055813 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X8 3 5 6 4 pmos1v_CDNS_7655933055814 $T=4560 -1510 0 0 $X=3880 $Y=-1710
X9 4 1 7 nmos1v_CDNS_7655933055815 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X10 3 2 6 4 pmos1v_CDNS_7655933055816 $T=1930 -1320 0 0 $X=1250 $Y=-1520
X11 3 6 1 4 pmos1v_CDNS_7655933055817 $T=2430 -1320 1 180 $X=1980 $Y=-1520
X12 6 2 7 4 nmos1v_CDNS_7655933055818 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y1 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=0
X0 1 M2_M1_CDNS_7655933055829 $T=80 250 0 0 $X=0 $Y=0
X1 2 M2_M1_CDNS_7655933055829 $T=480 250 0 0 $X=400 $Y=0
X2 3 M2_M1_CDNS_7655933055829 $T=880 250 0 0 $X=800 $Y=0
X3 4 M2_M1_CDNS_7655933055829 $T=1280 250 0 0 $X=1200 $Y=0
X4 5 M2_M1_CDNS_7655933055829 $T=1680 250 0 0 $X=1600 $Y=0
X5 6 M2_M1_CDNS_7655933055829 $T=2080 250 0 0 $X=2000 $Y=0
X6 7 M2_M1_CDNS_7655933055829 $T=2480 250 0 0 $X=2400 $Y=0
X7 8 M2_M1_CDNS_7655933055829 $T=2880 250 0 0 $X=2800 $Y=0
.ends MASCO__Y1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y2 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=0
X0 1 M3_M2_CDNS_765593305585 $T=80 250 0 0 $X=0 $Y=0
X1 2 M3_M2_CDNS_765593305585 $T=480 250 0 0 $X=400 $Y=0
X2 3 M3_M2_CDNS_765593305585 $T=880 250 0 0 $X=800 $Y=0
X3 4 M3_M2_CDNS_765593305585 $T=1280 250 0 0 $X=1200 $Y=0
X4 5 M3_M2_CDNS_765593305585 $T=1680 250 0 0 $X=1600 $Y=0
X5 6 M3_M2_CDNS_765593305585 $T=2080 250 0 0 $X=2000 $Y=0
X6 7 M3_M2_CDNS_765593305585 $T=2480 250 0 0 $X=2400 $Y=0
X7 8 M3_M2_CDNS_765593305585 $T=2880 250 0 0 $X=2800 $Y=0
.ends MASCO__Y2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceMultiplier                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceMultiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82
** N=210 EP=82 FDC=384
X0 1 M3_M2_CDNS_765593305585 $T=3380 31230 0 0 $X=3300 $Y=30980
X1 1 M3_M2_CDNS_765593305585 $T=3380 33140 0 0 $X=3300 $Y=32890
X2 1 M3_M2_CDNS_765593305585 $T=3380 34600 0 0 $X=3300 $Y=34350
X3 1 M3_M2_CDNS_765593305585 $T=3380 37680 0 0 $X=3300 $Y=37430
X4 1 M3_M2_CDNS_765593305585 $T=3380 39140 0 0 $X=3300 $Y=38890
X5 1 M3_M2_CDNS_765593305585 $T=3380 42220 0 0 $X=3300 $Y=41970
X6 1 M3_M2_CDNS_765593305585 $T=3380 43680 0 0 $X=3300 $Y=43430
X7 1 M3_M2_CDNS_765593305585 $T=3380 46750 0 0 $X=3300 $Y=46500
X8 1 M3_M2_CDNS_765593305585 $T=3380 48210 0 0 $X=3300 $Y=47960
X9 18 M3_M2_CDNS_765593305585 $T=8570 31230 0 0 $X=8490 $Y=30980
X10 18 M3_M2_CDNS_765593305585 $T=8570 33140 0 0 $X=8490 $Y=32890
X11 18 M3_M2_CDNS_765593305585 $T=8570 34600 0 0 $X=8490 $Y=34350
X12 18 M3_M2_CDNS_765593305585 $T=8570 37680 0 0 $X=8490 $Y=37430
X13 18 M3_M2_CDNS_765593305585 $T=8570 39140 0 0 $X=8490 $Y=38890
X14 18 M3_M2_CDNS_765593305585 $T=8570 42220 0 0 $X=8490 $Y=41970
X15 18 M3_M2_CDNS_765593305585 $T=8570 43680 0 0 $X=8490 $Y=43430
X16 18 M3_M2_CDNS_765593305585 $T=8570 46750 0 0 $X=8490 $Y=46500
X17 18 M3_M2_CDNS_765593305585 $T=8570 48210 0 0 $X=8490 $Y=47960
X18 26 M3_M2_CDNS_765593305585 $T=13600 31060 0 0 $X=13520 $Y=30810
X19 26 M3_M2_CDNS_765593305585 $T=13600 33140 0 0 $X=13520 $Y=32890
X20 26 M3_M2_CDNS_765593305585 $T=13600 34600 0 0 $X=13520 $Y=34350
X21 26 M3_M2_CDNS_765593305585 $T=13600 37680 0 0 $X=13520 $Y=37430
X22 26 M3_M2_CDNS_765593305585 $T=13600 39140 0 0 $X=13520 $Y=38890
X23 26 M3_M2_CDNS_765593305585 $T=13600 42220 0 0 $X=13520 $Y=41970
X24 26 M3_M2_CDNS_765593305585 $T=13600 43680 0 0 $X=13520 $Y=43430
X25 26 M3_M2_CDNS_765593305585 $T=13600 46750 0 0 $X=13520 $Y=46500
X26 26 M3_M2_CDNS_765593305585 $T=13600 48210 0 0 $X=13520 $Y=47960
X27 35 M3_M2_CDNS_765593305585 $T=18750 31230 0 0 $X=18670 $Y=30980
X28 35 M3_M2_CDNS_765593305585 $T=18750 33140 0 0 $X=18670 $Y=32890
X29 35 M3_M2_CDNS_765593305585 $T=18750 34600 0 0 $X=18670 $Y=34350
X30 35 M3_M2_CDNS_765593305585 $T=18750 37680 0 0 $X=18670 $Y=37430
X31 35 M3_M2_CDNS_765593305585 $T=18750 39140 0 0 $X=18670 $Y=38890
X32 35 M3_M2_CDNS_765593305585 $T=18750 42220 0 0 $X=18670 $Y=41970
X33 35 M3_M2_CDNS_765593305585 $T=18750 43680 0 0 $X=18670 $Y=43430
X34 35 M3_M2_CDNS_765593305585 $T=18750 46750 0 0 $X=18670 $Y=46500
X35 35 M3_M2_CDNS_765593305585 $T=18750 48210 0 0 $X=18670 $Y=47960
X36 44 M3_M2_CDNS_765593305585 $T=23840 31230 0 0 $X=23760 $Y=30980
X37 44 M3_M2_CDNS_765593305585 $T=23840 33140 0 0 $X=23760 $Y=32890
X38 44 M3_M2_CDNS_765593305585 $T=23840 34600 0 0 $X=23760 $Y=34350
X39 44 M3_M2_CDNS_765593305585 $T=23840 37680 0 0 $X=23760 $Y=37430
X40 44 M3_M2_CDNS_765593305585 $T=23840 39140 0 0 $X=23760 $Y=38890
X41 44 M3_M2_CDNS_765593305585 $T=23840 42220 0 0 $X=23760 $Y=41970
X42 44 M3_M2_CDNS_765593305585 $T=23840 43680 0 0 $X=23760 $Y=43430
X43 44 M3_M2_CDNS_765593305585 $T=23840 46750 0 0 $X=23760 $Y=46500
X44 44 M3_M2_CDNS_765593305585 $T=23840 48210 0 0 $X=23760 $Y=47960
X45 53 M3_M2_CDNS_765593305585 $T=28730 31230 0 0 $X=28650 $Y=30980
X46 53 M3_M2_CDNS_765593305585 $T=28730 33140 0 0 $X=28650 $Y=32890
X47 53 M3_M2_CDNS_765593305585 $T=28730 34600 0 0 $X=28650 $Y=34350
X48 53 M3_M2_CDNS_765593305585 $T=28730 37680 0 0 $X=28650 $Y=37430
X49 53 M3_M2_CDNS_765593305585 $T=28730 39140 0 0 $X=28650 $Y=38890
X50 53 M3_M2_CDNS_765593305585 $T=28730 42220 0 0 $X=28650 $Y=41970
X51 53 M3_M2_CDNS_765593305585 $T=28730 43680 0 0 $X=28650 $Y=43430
X52 53 M3_M2_CDNS_765593305585 $T=28730 46750 0 0 $X=28650 $Y=46500
X53 53 M3_M2_CDNS_765593305585 $T=28730 48210 0 0 $X=28650 $Y=47960
X54 62 M3_M2_CDNS_765593305585 $T=33970 31230 0 0 $X=33890 $Y=30980
X55 62 M3_M2_CDNS_765593305585 $T=33970 33140 0 0 $X=33890 $Y=32890
X56 62 M3_M2_CDNS_765593305585 $T=33970 34600 0 0 $X=33890 $Y=34350
X57 62 M3_M2_CDNS_765593305585 $T=33970 37680 0 0 $X=33890 $Y=37430
X58 62 M3_M2_CDNS_765593305585 $T=33970 39140 0 0 $X=33890 $Y=38890
X59 62 M3_M2_CDNS_765593305585 $T=33970 42220 0 0 $X=33890 $Y=41970
X60 62 M3_M2_CDNS_765593305585 $T=33970 43680 0 0 $X=33890 $Y=43430
X61 62 M3_M2_CDNS_765593305585 $T=33970 46750 0 0 $X=33890 $Y=46500
X62 62 M3_M2_CDNS_765593305585 $T=33970 48210 0 0 $X=33890 $Y=47960
X63 71 M3_M2_CDNS_765593305585 $T=39020 31230 0 0 $X=38940 $Y=30980
X64 71 M3_M2_CDNS_765593305585 $T=39020 33140 0 0 $X=38940 $Y=32890
X65 71 M3_M2_CDNS_765593305585 $T=39020 34600 0 0 $X=38940 $Y=34350
X66 71 M3_M2_CDNS_765593305585 $T=39020 37680 0 0 $X=38940 $Y=37430
X67 71 M3_M2_CDNS_765593305585 $T=39020 39140 0 0 $X=38940 $Y=38890
X68 71 M3_M2_CDNS_765593305585 $T=39020 42220 0 0 $X=38940 $Y=41970
X69 71 M3_M2_CDNS_765593305585 $T=39020 43680 0 0 $X=38940 $Y=43430
X70 71 M3_M2_CDNS_765593305585 $T=39020 46750 0 0 $X=38940 $Y=46500
X71 71 M3_M2_CDNS_765593305585 $T=39020 48210 0 0 $X=38940 $Y=47960
X72 2 M2_M1_CDNS_765593305586 $T=2220 31930 0 0 $X=2140 $Y=31800
X73 3 M2_M1_CDNS_765593305586 $T=2220 35820 0 0 $X=2140 $Y=35690
X74 4 M2_M1_CDNS_765593305586 $T=2220 36470 0 0 $X=2140 $Y=36340
X75 5 M2_M1_CDNS_765593305586 $T=2220 40360 0 0 $X=2140 $Y=40230
X76 6 M2_M1_CDNS_765593305586 $T=2220 41010 0 0 $X=2140 $Y=40880
X77 7 M2_M1_CDNS_765593305586 $T=2220 44900 0 0 $X=2140 $Y=44770
X78 8 M2_M1_CDNS_765593305586 $T=2220 45540 0 0 $X=2140 $Y=45410
X79 9 M2_M1_CDNS_765593305586 $T=2220 49430 0 0 $X=2140 $Y=49300
X80 2 M2_M1_CDNS_765593305586 $T=3380 32500 0 0 $X=3300 $Y=32370
X81 3 M2_M1_CDNS_765593305586 $T=3380 35240 0 0 $X=3300 $Y=35110
X82 4 M2_M1_CDNS_765593305586 $T=3380 37040 0 0 $X=3300 $Y=36910
X83 5 M2_M1_CDNS_765593305586 $T=3380 39780 0 0 $X=3300 $Y=39650
X84 6 M2_M1_CDNS_765593305586 $T=3380 41580 0 0 $X=3300 $Y=41450
X85 7 M2_M1_CDNS_765593305586 $T=3380 44320 0 0 $X=3300 $Y=44190
X86 8 M2_M1_CDNS_765593305586 $T=3380 46120 0 0 $X=3300 $Y=45990
X87 9 M2_M1_CDNS_765593305586 $T=3380 48860 0 0 $X=3300 $Y=48730
X88 2 M2_M1_CDNS_765593305586 $T=8590 32500 0 0 $X=8510 $Y=32370
X89 3 M2_M1_CDNS_765593305586 $T=8590 35240 0 0 $X=8510 $Y=35110
X90 4 M2_M1_CDNS_765593305586 $T=8590 37040 0 0 $X=8510 $Y=36910
X91 5 M2_M1_CDNS_765593305586 $T=8590 39780 0 0 $X=8510 $Y=39650
X92 6 M2_M1_CDNS_765593305586 $T=8590 41580 0 0 $X=8510 $Y=41450
X93 7 M2_M1_CDNS_765593305586 $T=8590 44320 0 0 $X=8510 $Y=44190
X94 8 M2_M1_CDNS_765593305586 $T=8590 46120 0 0 $X=8510 $Y=45990
X95 9 M2_M1_CDNS_765593305586 $T=8590 48860 0 0 $X=8510 $Y=48730
X96 2 M2_M1_CDNS_765593305586 $T=13610 32500 0 0 $X=13530 $Y=32370
X97 3 M2_M1_CDNS_765593305586 $T=13610 35240 0 0 $X=13530 $Y=35110
X98 4 M2_M1_CDNS_765593305586 $T=13610 37040 0 0 $X=13530 $Y=36910
X99 5 M2_M1_CDNS_765593305586 $T=13610 39780 0 0 $X=13530 $Y=39650
X100 6 M2_M1_CDNS_765593305586 $T=13610 41580 0 0 $X=13530 $Y=41450
X101 7 M2_M1_CDNS_765593305586 $T=13610 44320 0 0 $X=13530 $Y=44190
X102 8 M2_M1_CDNS_765593305586 $T=13610 46120 0 0 $X=13530 $Y=45990
X103 9 M2_M1_CDNS_765593305586 $T=13610 48860 0 0 $X=13530 $Y=48730
X104 2 M2_M1_CDNS_765593305586 $T=18740 32500 0 0 $X=18660 $Y=32370
X105 3 M2_M1_CDNS_765593305586 $T=18740 35240 0 0 $X=18660 $Y=35110
X106 4 M2_M1_CDNS_765593305586 $T=18740 37040 0 0 $X=18660 $Y=36910
X107 5 M2_M1_CDNS_765593305586 $T=18740 39780 0 0 $X=18660 $Y=39650
X108 6 M2_M1_CDNS_765593305586 $T=18740 41580 0 0 $X=18660 $Y=41450
X109 7 M2_M1_CDNS_765593305586 $T=18740 44320 0 0 $X=18660 $Y=44190
X110 8 M2_M1_CDNS_765593305586 $T=18740 46120 0 0 $X=18660 $Y=45990
X111 9 M2_M1_CDNS_765593305586 $T=18740 48860 0 0 $X=18660 $Y=48730
X112 2 M2_M1_CDNS_765593305586 $T=23810 32500 0 0 $X=23730 $Y=32370
X113 3 M2_M1_CDNS_765593305586 $T=23810 35240 0 0 $X=23730 $Y=35110
X114 4 M2_M1_CDNS_765593305586 $T=23810 37040 0 0 $X=23730 $Y=36910
X115 5 M2_M1_CDNS_765593305586 $T=23810 39780 0 0 $X=23730 $Y=39650
X116 6 M2_M1_CDNS_765593305586 $T=23810 41580 0 0 $X=23730 $Y=41450
X117 7 M2_M1_CDNS_765593305586 $T=23810 44320 0 0 $X=23730 $Y=44190
X118 8 M2_M1_CDNS_765593305586 $T=23810 46120 0 0 $X=23730 $Y=45990
X119 9 M2_M1_CDNS_765593305586 $T=23810 48860 0 0 $X=23730 $Y=48730
X120 2 M2_M1_CDNS_765593305586 $T=28690 32500 0 0 $X=28610 $Y=32370
X121 3 M2_M1_CDNS_765593305586 $T=28690 35240 0 0 $X=28610 $Y=35110
X122 4 M2_M1_CDNS_765593305586 $T=28690 37040 0 0 $X=28610 $Y=36910
X123 5 M2_M1_CDNS_765593305586 $T=28690 39780 0 0 $X=28610 $Y=39650
X124 6 M2_M1_CDNS_765593305586 $T=28690 41580 0 0 $X=28610 $Y=41450
X125 7 M2_M1_CDNS_765593305586 $T=28690 44320 0 0 $X=28610 $Y=44190
X126 8 M2_M1_CDNS_765593305586 $T=28690 46120 0 0 $X=28610 $Y=45990
X127 9 M2_M1_CDNS_765593305586 $T=28690 48860 0 0 $X=28610 $Y=48730
X128 2 M2_M1_CDNS_765593305586 $T=33890 32500 0 0 $X=33810 $Y=32370
X129 3 M2_M1_CDNS_765593305586 $T=33890 35240 0 0 $X=33810 $Y=35110
X130 4 M2_M1_CDNS_765593305586 $T=33890 37040 0 0 $X=33810 $Y=36910
X131 5 M2_M1_CDNS_765593305586 $T=33890 39780 0 0 $X=33810 $Y=39650
X132 6 M2_M1_CDNS_765593305586 $T=33890 41580 0 0 $X=33810 $Y=41450
X133 7 M2_M1_CDNS_765593305586 $T=33890 44320 0 0 $X=33810 $Y=44190
X134 8 M2_M1_CDNS_765593305586 $T=33890 46120 0 0 $X=33810 $Y=45990
X135 9 M2_M1_CDNS_765593305586 $T=33890 48860 0 0 $X=33810 $Y=48730
X136 2 M2_M1_CDNS_765593305586 $T=38920 32500 0 0 $X=38840 $Y=32370
X137 3 M2_M1_CDNS_765593305586 $T=38920 35240 0 0 $X=38840 $Y=35110
X138 4 M2_M1_CDNS_765593305586 $T=38920 37040 0 0 $X=38840 $Y=36910
X139 5 M2_M1_CDNS_765593305586 $T=38920 39780 0 0 $X=38840 $Y=39650
X140 6 M2_M1_CDNS_765593305586 $T=38920 41580 0 0 $X=38840 $Y=41450
X141 7 M2_M1_CDNS_765593305586 $T=38920 44320 0 0 $X=38840 $Y=44190
X142 8 M2_M1_CDNS_765593305586 $T=38920 46120 0 0 $X=38840 $Y=45990
X143 9 M2_M1_CDNS_765593305586 $T=38920 48860 0 0 $X=38840 $Y=48730
X144 1 M2_M1_CDNS_7655933055829 $T=3380 31230 0 0 $X=3300 $Y=30980
X145 1 M2_M1_CDNS_7655933055829 $T=3380 33140 0 0 $X=3300 $Y=32890
X146 1 M2_M1_CDNS_7655933055829 $T=3380 34600 0 0 $X=3300 $Y=34350
X147 1 M2_M1_CDNS_7655933055829 $T=3380 37680 0 0 $X=3300 $Y=37430
X148 1 M2_M1_CDNS_7655933055829 $T=3380 39140 0 0 $X=3300 $Y=38890
X149 1 M2_M1_CDNS_7655933055829 $T=3380 42220 0 0 $X=3300 $Y=41970
X150 1 M2_M1_CDNS_7655933055829 $T=3380 43680 0 0 $X=3300 $Y=43430
X151 1 M2_M1_CDNS_7655933055829 $T=3380 46750 0 0 $X=3300 $Y=46500
X152 1 M2_M1_CDNS_7655933055829 $T=3380 48210 0 0 $X=3300 $Y=47960
X153 18 M2_M1_CDNS_7655933055829 $T=8570 31230 0 0 $X=8490 $Y=30980
X154 18 M2_M1_CDNS_7655933055829 $T=8570 33140 0 0 $X=8490 $Y=32890
X155 18 M2_M1_CDNS_7655933055829 $T=8570 34600 0 0 $X=8490 $Y=34350
X156 18 M2_M1_CDNS_7655933055829 $T=8570 37680 0 0 $X=8490 $Y=37430
X157 18 M2_M1_CDNS_7655933055829 $T=8570 39140 0 0 $X=8490 $Y=38890
X158 18 M2_M1_CDNS_7655933055829 $T=8570 42220 0 0 $X=8490 $Y=41970
X159 18 M2_M1_CDNS_7655933055829 $T=8570 43680 0 0 $X=8490 $Y=43430
X160 18 M2_M1_CDNS_7655933055829 $T=8570 46750 0 0 $X=8490 $Y=46500
X161 18 M2_M1_CDNS_7655933055829 $T=8570 48210 0 0 $X=8490 $Y=47960
X162 26 M2_M1_CDNS_7655933055829 $T=13600 31060 0 0 $X=13520 $Y=30810
X163 26 M2_M1_CDNS_7655933055829 $T=13600 33140 0 0 $X=13520 $Y=32890
X164 26 M2_M1_CDNS_7655933055829 $T=13600 34600 0 0 $X=13520 $Y=34350
X165 26 M2_M1_CDNS_7655933055829 $T=13600 37680 0 0 $X=13520 $Y=37430
X166 26 M2_M1_CDNS_7655933055829 $T=13600 39140 0 0 $X=13520 $Y=38890
X167 26 M2_M1_CDNS_7655933055829 $T=13600 42220 0 0 $X=13520 $Y=41970
X168 26 M2_M1_CDNS_7655933055829 $T=13600 43680 0 0 $X=13520 $Y=43430
X169 26 M2_M1_CDNS_7655933055829 $T=13600 46750 0 0 $X=13520 $Y=46500
X170 26 M2_M1_CDNS_7655933055829 $T=13600 48210 0 0 $X=13520 $Y=47960
X171 35 M2_M1_CDNS_7655933055829 $T=18750 31230 0 0 $X=18670 $Y=30980
X172 35 M2_M1_CDNS_7655933055829 $T=18750 33140 0 0 $X=18670 $Y=32890
X173 35 M2_M1_CDNS_7655933055829 $T=18750 34600 0 0 $X=18670 $Y=34350
X174 35 M2_M1_CDNS_7655933055829 $T=18750 37680 0 0 $X=18670 $Y=37430
X175 35 M2_M1_CDNS_7655933055829 $T=18750 39140 0 0 $X=18670 $Y=38890
X176 35 M2_M1_CDNS_7655933055829 $T=18750 42220 0 0 $X=18670 $Y=41970
X177 35 M2_M1_CDNS_7655933055829 $T=18750 43680 0 0 $X=18670 $Y=43430
X178 35 M2_M1_CDNS_7655933055829 $T=18750 46750 0 0 $X=18670 $Y=46500
X179 35 M2_M1_CDNS_7655933055829 $T=18750 48210 0 0 $X=18670 $Y=47960
X180 44 M2_M1_CDNS_7655933055829 $T=23840 31230 0 0 $X=23760 $Y=30980
X181 44 M2_M1_CDNS_7655933055829 $T=23840 33140 0 0 $X=23760 $Y=32890
X182 44 M2_M1_CDNS_7655933055829 $T=23840 34600 0 0 $X=23760 $Y=34350
X183 44 M2_M1_CDNS_7655933055829 $T=23840 37680 0 0 $X=23760 $Y=37430
X184 44 M2_M1_CDNS_7655933055829 $T=23840 39140 0 0 $X=23760 $Y=38890
X185 44 M2_M1_CDNS_7655933055829 $T=23840 42220 0 0 $X=23760 $Y=41970
X186 44 M2_M1_CDNS_7655933055829 $T=23840 43680 0 0 $X=23760 $Y=43430
X187 44 M2_M1_CDNS_7655933055829 $T=23840 46750 0 0 $X=23760 $Y=46500
X188 44 M2_M1_CDNS_7655933055829 $T=23840 48210 0 0 $X=23760 $Y=47960
X189 53 M2_M1_CDNS_7655933055829 $T=28730 31230 0 0 $X=28650 $Y=30980
X190 53 M2_M1_CDNS_7655933055829 $T=28730 33140 0 0 $X=28650 $Y=32890
X191 53 M2_M1_CDNS_7655933055829 $T=28730 34600 0 0 $X=28650 $Y=34350
X192 53 M2_M1_CDNS_7655933055829 $T=28730 37680 0 0 $X=28650 $Y=37430
X193 53 M2_M1_CDNS_7655933055829 $T=28730 39140 0 0 $X=28650 $Y=38890
X194 53 M2_M1_CDNS_7655933055829 $T=28730 42220 0 0 $X=28650 $Y=41970
X195 53 M2_M1_CDNS_7655933055829 $T=28730 43680 0 0 $X=28650 $Y=43430
X196 53 M2_M1_CDNS_7655933055829 $T=28730 46750 0 0 $X=28650 $Y=46500
X197 53 M2_M1_CDNS_7655933055829 $T=28730 48210 0 0 $X=28650 $Y=47960
X198 62 M2_M1_CDNS_7655933055829 $T=33970 31230 0 0 $X=33890 $Y=30980
X199 62 M2_M1_CDNS_7655933055829 $T=33970 33140 0 0 $X=33890 $Y=32890
X200 62 M2_M1_CDNS_7655933055829 $T=33970 34600 0 0 $X=33890 $Y=34350
X201 62 M2_M1_CDNS_7655933055829 $T=33970 37680 0 0 $X=33890 $Y=37430
X202 62 M2_M1_CDNS_7655933055829 $T=33970 39140 0 0 $X=33890 $Y=38890
X203 62 M2_M1_CDNS_7655933055829 $T=33970 42220 0 0 $X=33890 $Y=41970
X204 62 M2_M1_CDNS_7655933055829 $T=33970 43680 0 0 $X=33890 $Y=43430
X205 62 M2_M1_CDNS_7655933055829 $T=33970 46750 0 0 $X=33890 $Y=46500
X206 62 M2_M1_CDNS_7655933055829 $T=33970 48210 0 0 $X=33890 $Y=47960
X207 71 M2_M1_CDNS_7655933055829 $T=39020 31230 0 0 $X=38940 $Y=30980
X208 71 M2_M1_CDNS_7655933055829 $T=39020 33140 0 0 $X=38940 $Y=32890
X209 71 M2_M1_CDNS_7655933055829 $T=39020 34600 0 0 $X=38940 $Y=34350
X210 71 M2_M1_CDNS_7655933055829 $T=39020 37680 0 0 $X=38940 $Y=37430
X211 71 M2_M1_CDNS_7655933055829 $T=39020 39140 0 0 $X=38940 $Y=38890
X212 71 M2_M1_CDNS_7655933055829 $T=39020 42220 0 0 $X=38940 $Y=41970
X213 71 M2_M1_CDNS_7655933055829 $T=39020 43680 0 0 $X=38940 $Y=43430
X214 71 M2_M1_CDNS_7655933055829 $T=39020 46750 0 0 $X=38940 $Y=46500
X215 71 M2_M1_CDNS_7655933055829 $T=39020 48210 0 0 $X=38940 $Y=47960
X216 1 2 10 11 19 90 154 AND $T=2730 30830 1 0 $X=3800 $Y=31540
X217 1 3 10 11 20 89 153 AND $T=2730 36910 0 0 $X=3800 $Y=33810
X218 1 4 10 11 12 88 152 AND $T=2730 35370 1 0 $X=3800 $Y=36080
X219 1 5 10 11 13 87 151 AND $T=2730 41450 0 0 $X=3800 $Y=38350
X220 1 6 10 11 14 86 150 AND $T=2730 39910 1 0 $X=3800 $Y=40620
X221 1 7 10 11 15 85 149 AND $T=2730 45990 0 0 $X=3800 $Y=42890
X222 1 8 10 11 16 84 148 AND $T=2730 44450 1 0 $X=3800 $Y=45160
X223 1 9 10 11 17 83 147 AND $T=2730 50530 0 0 $X=3800 $Y=47430
X224 18 2 10 11 27 98 162 AND $T=7940 30820 1 0 $X=9010 $Y=31530
X225 18 3 10 11 28 97 161 AND $T=7940 36900 0 0 $X=9010 $Y=33800
X226 18 4 10 11 29 96 160 AND $T=7940 35370 1 0 $X=9010 $Y=36080
X227 18 5 10 11 21 95 159 AND $T=7940 41450 0 0 $X=9010 $Y=38350
X228 18 6 10 11 22 94 158 AND $T=7940 39910 1 0 $X=9010 $Y=40620
X229 18 7 10 11 23 93 157 AND $T=7940 45990 0 0 $X=9010 $Y=42890
X230 18 8 10 11 24 92 156 AND $T=7940 44450 1 0 $X=9010 $Y=45160
X231 18 9 10 11 25 91 155 AND $T=7940 50530 0 0 $X=9010 $Y=47430
X232 26 2 10 11 36 106 170 AND $T=12940 30820 1 0 $X=14010 $Y=31530
X233 26 3 10 11 37 105 169 AND $T=12940 36900 0 0 $X=14010 $Y=33800
X234 26 4 10 11 38 104 168 AND $T=12940 35370 1 0 $X=14010 $Y=36080
X235 26 5 10 11 30 103 167 AND $T=12940 41450 0 0 $X=14010 $Y=38350
X236 26 6 10 11 31 102 166 AND $T=12940 39910 1 0 $X=14010 $Y=40620
X237 26 7 10 11 32 101 165 AND $T=12940 45990 0 0 $X=14010 $Y=42890
X238 26 8 10 11 33 100 164 AND $T=12940 44450 1 0 $X=14010 $Y=45160
X239 26 9 10 11 34 99 163 AND $T=12940 50530 0 0 $X=14010 $Y=47430
X240 35 2 10 11 45 114 178 AND $T=18070 30820 1 0 $X=19140 $Y=31530
X241 35 3 10 11 46 113 177 AND $T=18070 36900 0 0 $X=19140 $Y=33800
X242 35 4 10 11 47 112 176 AND $T=18070 35370 1 0 $X=19140 $Y=36080
X243 35 5 10 11 39 111 175 AND $T=18070 41450 0 0 $X=19140 $Y=38350
X244 35 6 10 11 40 110 174 AND $T=18070 39910 1 0 $X=19140 $Y=40620
X245 35 7 10 11 41 109 173 AND $T=18070 45990 0 0 $X=19140 $Y=42890
X246 35 8 10 11 42 108 172 AND $T=18070 44450 1 0 $X=19140 $Y=45160
X247 35 9 10 11 43 107 171 AND $T=18070 50530 0 0 $X=19140 $Y=47430
X248 44 2 10 11 54 122 186 AND $T=23140 30820 1 0 $X=24210 $Y=31530
X249 44 3 10 11 55 121 185 AND $T=23140 36900 0 0 $X=24210 $Y=33800
X250 44 4 10 11 56 120 184 AND $T=23140 35370 1 0 $X=24210 $Y=36080
X251 44 5 10 11 48 119 183 AND $T=23140 41450 0 0 $X=24210 $Y=38350
X252 44 6 10 11 49 118 182 AND $T=23140 39910 1 0 $X=24210 $Y=40620
X253 44 7 10 11 50 117 181 AND $T=23140 45990 0 0 $X=24210 $Y=42890
X254 44 8 10 11 51 116 180 AND $T=23140 44450 1 0 $X=24210 $Y=45160
X255 44 9 10 11 52 115 179 AND $T=23140 50530 0 0 $X=24210 $Y=47430
X256 53 2 10 11 63 130 194 AND $T=28010 30820 1 0 $X=29080 $Y=31530
X257 53 3 10 11 64 129 193 AND $T=28010 36900 0 0 $X=29080 $Y=33800
X258 53 4 10 11 65 128 192 AND $T=28010 35370 1 0 $X=29080 $Y=36080
X259 53 5 10 11 57 127 191 AND $T=28010 41450 0 0 $X=29080 $Y=38350
X260 53 6 10 11 58 126 190 AND $T=28010 39910 1 0 $X=29080 $Y=40620
X261 53 7 10 11 59 125 189 AND $T=28010 45990 0 0 $X=29080 $Y=42890
X262 53 8 10 11 60 124 188 AND $T=28010 44450 1 0 $X=29080 $Y=45160
X263 53 9 10 11 61 123 187 AND $T=28010 50530 0 0 $X=29080 $Y=47430
X264 62 2 10 11 72 138 202 AND $T=33230 30830 1 0 $X=34300 $Y=31540
X265 62 3 10 11 73 137 201 AND $T=33230 36900 0 0 $X=34300 $Y=33800
X266 62 4 10 11 74 136 200 AND $T=33230 35370 1 0 $X=34300 $Y=36080
X267 62 5 10 11 66 135 199 AND $T=33230 41450 0 0 $X=34300 $Y=38350
X268 62 6 10 11 67 134 198 AND $T=33230 39910 1 0 $X=34300 $Y=40620
X269 62 7 10 11 68 133 197 AND $T=33230 45990 0 0 $X=34300 $Y=42890
X270 62 8 10 11 69 132 196 AND $T=33230 44450 1 0 $X=34300 $Y=45160
X271 62 9 10 11 70 131 195 AND $T=33230 50530 0 0 $X=34300 $Y=47430
X272 71 2 10 11 80 146 210 AND $T=38250 30830 1 0 $X=39320 $Y=31540
X273 71 3 10 11 81 145 209 AND $T=38250 36910 0 0 $X=39320 $Y=33810
X274 71 4 10 11 82 144 208 AND $T=38250 35370 1 0 $X=39320 $Y=36080
X275 71 5 10 11 75 143 207 AND $T=38250 41450 0 0 $X=39320 $Y=38350
X276 71 6 10 11 76 142 206 AND $T=38250 39910 1 0 $X=39320 $Y=40620
X277 71 7 10 11 77 141 205 AND $T=38250 45990 0 0 $X=39320 $Y=42890
X278 71 8 10 11 78 140 204 AND $T=38250 44450 1 0 $X=39320 $Y=45160
X279 71 9 10 11 79 139 203 AND $T=38250 50530 0 0 $X=39320 $Y=47430
X280 17 16 15 14 13 12 20 19 MASCO__Y1 $T=4320 31030 0 0 $X=4320 $Y=31030
X281 25 24 23 22 21 29 28 27 MASCO__Y1 $T=9530 31030 0 0 $X=9530 $Y=31030
X282 34 33 32 31 30 38 37 36 MASCO__Y1 $T=14515 31030 0 0 $X=14515 $Y=31030
X283 43 42 41 40 39 47 46 45 MASCO__Y1 $T=19655 31030 0 0 $X=19655 $Y=31030
X284 52 51 50 49 48 56 55 54 MASCO__Y1 $T=24735 31030 0 0 $X=24735 $Y=31030
X285 61 60 59 58 57 65 64 63 MASCO__Y1 $T=29595 31030 0 0 $X=29595 $Y=31030
X286 70 69 68 67 66 74 73 72 MASCO__Y1 $T=34815 31030 0 0 $X=34815 $Y=31030
X287 79 78 77 76 75 82 81 80 MASCO__Y1 $T=39840 31030 0 0 $X=39840 $Y=31030
X288 17 16 15 14 13 12 20 19 MASCO__Y2 $T=4320 31030 0 0 $X=4320 $Y=31030
X289 25 24 23 22 21 29 28 27 MASCO__Y2 $T=9530 31030 0 0 $X=9530 $Y=31030
X290 34 33 32 31 30 38 37 36 MASCO__Y2 $T=14515 31030 0 0 $X=14515 $Y=31030
X291 43 42 41 40 39 47 46 45 MASCO__Y2 $T=19655 31030 0 0 $X=19655 $Y=31030
X292 52 51 50 49 48 56 55 54 MASCO__Y2 $T=24735 31030 0 0 $X=24735 $Y=31030
X293 61 60 59 58 57 65 64 63 MASCO__Y2 $T=29595 31030 0 0 $X=29595 $Y=31030
X294 70 69 68 67 66 74 73 72 MASCO__Y2 $T=34815 31030 0 0 $X=34815 $Y=31030
X295 79 78 77 76 75 82 81 80 MASCO__Y2 $T=39840 31030 0 0 $X=39840 $Y=31030
M0 154 2 90 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=33350 $dt=0
M1 153 3 89 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=34150 $dt=0
M2 152 4 88 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=37890 $dt=0
M3 151 5 87 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=38690 $dt=0
M4 150 6 86 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=42430 $dt=0
M5 149 7 85 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=43230 $dt=0
M6 148 8 84 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=46970 $dt=0
M7 147 9 83 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=47770 $dt=0
M8 11 1 154 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=33350 $dt=0
M9 11 1 153 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=34150 $dt=0
M10 11 1 152 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=37890 $dt=0
M11 11 1 151 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=38690 $dt=0
M12 11 1 150 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=42430 $dt=0
M13 11 1 149 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=43230 $dt=0
M14 11 1 148 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=46970 $dt=0
M15 11 1 147 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=47770 $dt=0
M16 19 90 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=33360 $dt=0
M17 20 89 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=34140 $dt=0
M18 12 88 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=37900 $dt=0
M19 13 87 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=38680 $dt=0
M20 14 86 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=42440 $dt=0
M21 15 85 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=43220 $dt=0
M22 16 84 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=46980 $dt=0
M23 17 83 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=47760 $dt=0
M24 162 2 98 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=33340 $dt=0
M25 161 3 97 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=34140 $dt=0
M26 160 4 96 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=37890 $dt=0
M27 159 5 95 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=38690 $dt=0
M28 158 6 94 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=42430 $dt=0
M29 157 7 93 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=43230 $dt=0
M30 156 8 92 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=46970 $dt=0
M31 155 9 91 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=47770 $dt=0
M32 11 18 162 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=33340 $dt=0
M33 11 18 161 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=34140 $dt=0
M34 11 18 160 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=37890 $dt=0
M35 11 18 159 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=38690 $dt=0
M36 11 18 158 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=42430 $dt=0
M37 11 18 157 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=43230 $dt=0
M38 11 18 156 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=46970 $dt=0
M39 11 18 155 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=47770 $dt=0
M40 27 98 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=33350 $dt=0
M41 28 97 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=34130 $dt=0
M42 29 96 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=37900 $dt=0
M43 21 95 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=38680 $dt=0
M44 22 94 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=42440 $dt=0
M45 23 93 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=43220 $dt=0
M46 24 92 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=46980 $dt=0
M47 25 91 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=47760 $dt=0
M48 170 2 106 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=33340 $dt=0
M49 169 3 105 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=34140 $dt=0
M50 168 4 104 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=37890 $dt=0
M51 167 5 103 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=38690 $dt=0
M52 166 6 102 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=42430 $dt=0
M53 165 7 101 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=43230 $dt=0
M54 164 8 100 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=46970 $dt=0
M55 163 9 99 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=47770 $dt=0
M56 11 26 170 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=33340 $dt=0
M57 11 26 169 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=34140 $dt=0
M58 11 26 168 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=37890 $dt=0
M59 11 26 167 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=38690 $dt=0
M60 11 26 166 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=42430 $dt=0
M61 11 26 165 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=43230 $dt=0
M62 11 26 164 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=46970 $dt=0
M63 11 26 163 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=47770 $dt=0
M64 36 106 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=33350 $dt=0
M65 37 105 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=34130 $dt=0
M66 38 104 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=37900 $dt=0
M67 30 103 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=38680 $dt=0
M68 31 102 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=42440 $dt=0
M69 32 101 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=43220 $dt=0
M70 33 100 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=46980 $dt=0
M71 34 99 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=47760 $dt=0
M72 178 2 114 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=33340 $dt=0
M73 177 3 113 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=34140 $dt=0
M74 176 4 112 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=37890 $dt=0
M75 175 5 111 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=38690 $dt=0
M76 174 6 110 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=42430 $dt=0
M77 173 7 109 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=43230 $dt=0
M78 172 8 108 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=46970 $dt=0
M79 171 9 107 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=47770 $dt=0
M80 11 35 178 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=33340 $dt=0
M81 11 35 177 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=34140 $dt=0
M82 11 35 176 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=37890 $dt=0
M83 11 35 175 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=38690 $dt=0
M84 11 35 174 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=42430 $dt=0
M85 11 35 173 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=43230 $dt=0
M86 11 35 172 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=46970 $dt=0
M87 11 35 171 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=47770 $dt=0
M88 45 114 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=33350 $dt=0
M89 46 113 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=34130 $dt=0
M90 47 112 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=37900 $dt=0
M91 39 111 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=38680 $dt=0
M92 40 110 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=42440 $dt=0
M93 41 109 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=43220 $dt=0
M94 42 108 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=46980 $dt=0
M95 43 107 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=47760 $dt=0
M96 186 2 122 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=33340 $dt=0
M97 185 3 121 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=34140 $dt=0
M98 184 4 120 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=37890 $dt=0
M99 183 5 119 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=38690 $dt=0
M100 182 6 118 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=42430 $dt=0
M101 181 7 117 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=43230 $dt=0
M102 180 8 116 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=46970 $dt=0
M103 179 9 115 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=47770 $dt=0
M104 11 44 186 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=33340 $dt=0
M105 11 44 185 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=34140 $dt=0
M106 11 44 184 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=37890 $dt=0
M107 11 44 183 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=38690 $dt=0
M108 11 44 182 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=42430 $dt=0
M109 11 44 181 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=43230 $dt=0
M110 11 44 180 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=46970 $dt=0
M111 11 44 179 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=47770 $dt=0
M112 54 122 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=33350 $dt=0
M113 55 121 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=34130 $dt=0
M114 56 120 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=37900 $dt=0
M115 48 119 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=38680 $dt=0
M116 49 118 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=42440 $dt=0
M117 50 117 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=43220 $dt=0
M118 51 116 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=46980 $dt=0
M119 52 115 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=47760 $dt=0
M120 194 2 130 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=33340 $dt=0
M121 193 3 129 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=34140 $dt=0
M122 192 4 128 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=37890 $dt=0
M123 191 5 127 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=38690 $dt=0
M124 190 6 126 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=42430 $dt=0
M125 189 7 125 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=43230 $dt=0
M126 188 8 124 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=46970 $dt=0
M127 187 9 123 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=47770 $dt=0
M128 11 53 194 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=33340 $dt=0
M129 11 53 193 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=34140 $dt=0
M130 11 53 192 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=37890 $dt=0
M131 11 53 191 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=38690 $dt=0
M132 11 53 190 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=42430 $dt=0
M133 11 53 189 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=43230 $dt=0
M134 11 53 188 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=46970 $dt=0
M135 11 53 187 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=47770 $dt=0
M136 63 130 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=33350 $dt=0
M137 64 129 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=34130 $dt=0
M138 65 128 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=37900 $dt=0
M139 57 127 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=38680 $dt=0
M140 58 126 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=42440 $dt=0
M141 59 125 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=43220 $dt=0
M142 60 124 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=46980 $dt=0
M143 61 123 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=47760 $dt=0
M144 202 2 138 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=33350 $dt=0
M145 201 3 137 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=34140 $dt=0
M146 200 4 136 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=37890 $dt=0
M147 199 5 135 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=38690 $dt=0
M148 198 6 134 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=42430 $dt=0
M149 197 7 133 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=43230 $dt=0
M150 196 8 132 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=46970 $dt=0
M151 195 9 131 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=47770 $dt=0
M152 11 62 202 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=33350 $dt=0
M153 11 62 201 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=34140 $dt=0
M154 11 62 200 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=37890 $dt=0
M155 11 62 199 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=38690 $dt=0
M156 11 62 198 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=42430 $dt=0
M157 11 62 197 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=43230 $dt=0
M158 11 62 196 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=46970 $dt=0
M159 11 62 195 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=47770 $dt=0
M160 72 138 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=33360 $dt=0
M161 73 137 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=34130 $dt=0
M162 74 136 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=37900 $dt=0
M163 66 135 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=38680 $dt=0
M164 67 134 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=42440 $dt=0
M165 68 133 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=43220 $dt=0
M166 69 132 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=46980 $dt=0
M167 70 131 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=47760 $dt=0
M168 210 2 146 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=33350 $dt=0
M169 209 3 145 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=34150 $dt=0
M170 208 4 144 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=37890 $dt=0
M171 207 5 143 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=38690 $dt=0
M172 206 6 142 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=42430 $dt=0
M173 205 7 141 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=43230 $dt=0
M174 204 8 140 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=46970 $dt=0
M175 203 9 139 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=47770 $dt=0
M176 11 71 210 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=33350 $dt=0
M177 11 71 209 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=34150 $dt=0
M178 11 71 208 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=37890 $dt=0
M179 11 71 207 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=38690 $dt=0
M180 11 71 206 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=42430 $dt=0
M181 11 71 205 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=43230 $dt=0
M182 11 71 204 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=46970 $dt=0
M183 11 71 203 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=47770 $dt=0
M184 80 146 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=33360 $dt=0
M185 81 145 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=34140 $dt=0
M186 82 144 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=37900 $dt=0
M187 75 143 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=38680 $dt=0
M188 76 142 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=42440 $dt=0
M189 77 141 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=43220 $dt=0
M190 78 140 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=46980 $dt=0
M191 79 139 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=47760 $dt=0
M192 90 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=31910 $dt=1
M193 89 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=35590 $dt=1
M194 88 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=36450 $dt=1
M195 87 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40130 $dt=1
M196 86 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40990 $dt=1
M197 85 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=44670 $dt=1
M198 84 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=45530 $dt=1
M199 83 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=49210 $dt=1
M200 10 1 90 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=31910 $dt=1
M201 10 1 89 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=35590 $dt=1
M202 10 1 88 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=36450 $dt=1
M203 10 1 87 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40130 $dt=1
M204 10 1 86 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40990 $dt=1
M205 10 1 85 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=44670 $dt=1
M206 10 1 84 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=45530 $dt=1
M207 10 1 83 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=49210 $dt=1
M208 19 90 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=31860 $dt=1
M209 20 89 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=35400 $dt=1
M210 12 88 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=36400 $dt=1
M211 13 87 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=39940 $dt=1
M212 14 86 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=40940 $dt=1
M213 15 85 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=44480 $dt=1
M214 16 84 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=45480 $dt=1
M215 17 83 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=49020 $dt=1
M216 98 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=31900 $dt=1
M217 97 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=35580 $dt=1
M218 96 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=36450 $dt=1
M219 95 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40130 $dt=1
M220 94 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40990 $dt=1
M221 93 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=44670 $dt=1
M222 92 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=45530 $dt=1
M223 91 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=49210 $dt=1
M224 10 18 98 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=31900 $dt=1
M225 10 18 97 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=35580 $dt=1
M226 10 18 96 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=36450 $dt=1
M227 10 18 95 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40130 $dt=1
M228 10 18 94 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40990 $dt=1
M229 10 18 93 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=44670 $dt=1
M230 10 18 92 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=45530 $dt=1
M231 10 18 91 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=49210 $dt=1
M232 27 98 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=31850 $dt=1
M233 28 97 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=35390 $dt=1
M234 29 96 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=36400 $dt=1
M235 21 95 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=39940 $dt=1
M236 22 94 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=40940 $dt=1
M237 23 93 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=44480 $dt=1
M238 24 92 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=45480 $dt=1
M239 25 91 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=49020 $dt=1
M240 106 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=31900 $dt=1
M241 105 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=35580 $dt=1
M242 104 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=36450 $dt=1
M243 103 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40130 $dt=1
M244 102 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40990 $dt=1
M245 101 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=44670 $dt=1
M246 100 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=45530 $dt=1
M247 99 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=49210 $dt=1
M248 10 26 106 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=31900 $dt=1
M249 10 26 105 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=35580 $dt=1
M250 10 26 104 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=36450 $dt=1
M251 10 26 103 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40130 $dt=1
M252 10 26 102 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40990 $dt=1
M253 10 26 101 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=44670 $dt=1
M254 10 26 100 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=45530 $dt=1
M255 10 26 99 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=49210 $dt=1
M256 36 106 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=31850 $dt=1
M257 37 105 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=35390 $dt=1
M258 38 104 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=36400 $dt=1
M259 30 103 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=39940 $dt=1
M260 31 102 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=40940 $dt=1
M261 32 101 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=44480 $dt=1
M262 33 100 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=45480 $dt=1
M263 34 99 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=49020 $dt=1
M264 114 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=31900 $dt=1
M265 113 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=35580 $dt=1
M266 112 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=36450 $dt=1
M267 111 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40130 $dt=1
M268 110 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40990 $dt=1
M269 109 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=44670 $dt=1
M270 108 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=45530 $dt=1
M271 107 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=49210 $dt=1
M272 10 35 114 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=31900 $dt=1
M273 10 35 113 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=35580 $dt=1
M274 10 35 112 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=36450 $dt=1
M275 10 35 111 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40130 $dt=1
M276 10 35 110 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40990 $dt=1
M277 10 35 109 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=44670 $dt=1
M278 10 35 108 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=45530 $dt=1
M279 10 35 107 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=49210 $dt=1
M280 45 114 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=31850 $dt=1
M281 46 113 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=35390 $dt=1
M282 47 112 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=36400 $dt=1
M283 39 111 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=39940 $dt=1
M284 40 110 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=40940 $dt=1
M285 41 109 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=44480 $dt=1
M286 42 108 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=45480 $dt=1
M287 43 107 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=49020 $dt=1
M288 122 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=31900 $dt=1
M289 121 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=35580 $dt=1
M290 120 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=36450 $dt=1
M291 119 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40130 $dt=1
M292 118 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40990 $dt=1
M293 117 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=44670 $dt=1
M294 116 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=45530 $dt=1
M295 115 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=49210 $dt=1
M296 10 44 122 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=31900 $dt=1
M297 10 44 121 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=35580 $dt=1
M298 10 44 120 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=36450 $dt=1
M299 10 44 119 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40130 $dt=1
M300 10 44 118 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40990 $dt=1
M301 10 44 117 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=44670 $dt=1
M302 10 44 116 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=45530 $dt=1
M303 10 44 115 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=49210 $dt=1
M304 54 122 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=31850 $dt=1
M305 55 121 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=35390 $dt=1
M306 56 120 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=36400 $dt=1
M307 48 119 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=39940 $dt=1
M308 49 118 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=40940 $dt=1
M309 50 117 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=44480 $dt=1
M310 51 116 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=45480 $dt=1
M311 52 115 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=49020 $dt=1
M312 130 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=31900 $dt=1
M313 129 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=35580 $dt=1
M314 128 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=36450 $dt=1
M315 127 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40130 $dt=1
M316 126 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40990 $dt=1
M317 125 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=44670 $dt=1
M318 124 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=45530 $dt=1
M319 123 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=49210 $dt=1
M320 10 53 130 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=31900 $dt=1
M321 10 53 129 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=35580 $dt=1
M322 10 53 128 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=36450 $dt=1
M323 10 53 127 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40130 $dt=1
M324 10 53 126 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40990 $dt=1
M325 10 53 125 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=44670 $dt=1
M326 10 53 124 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=45530 $dt=1
M327 10 53 123 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=49210 $dt=1
M328 63 130 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=31850 $dt=1
M329 64 129 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=35390 $dt=1
M330 65 128 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=36400 $dt=1
M331 57 127 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=39940 $dt=1
M332 58 126 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=40940 $dt=1
M333 59 125 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=44480 $dt=1
M334 60 124 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=45480 $dt=1
M335 61 123 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=49020 $dt=1
M336 138 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=31910 $dt=1
M337 137 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=35580 $dt=1
M338 136 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=36450 $dt=1
M339 135 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40130 $dt=1
M340 134 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40990 $dt=1
M341 133 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=44670 $dt=1
M342 132 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=45530 $dt=1
M343 131 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=49210 $dt=1
M344 10 62 138 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=31910 $dt=1
M345 10 62 137 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=35580 $dt=1
M346 10 62 136 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=36450 $dt=1
M347 10 62 135 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40130 $dt=1
M348 10 62 134 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40990 $dt=1
M349 10 62 133 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=44670 $dt=1
M350 10 62 132 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=45530 $dt=1
M351 10 62 131 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=49210 $dt=1
M352 72 138 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=31860 $dt=1
M353 73 137 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=35390 $dt=1
M354 74 136 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=36400 $dt=1
M355 66 135 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=39940 $dt=1
M356 67 134 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=40940 $dt=1
M357 68 133 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=44480 $dt=1
M358 69 132 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=45480 $dt=1
M359 70 131 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=49020 $dt=1
M360 146 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=31910 $dt=1
M361 145 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=35590 $dt=1
M362 144 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=36450 $dt=1
M363 143 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40130 $dt=1
M364 142 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40990 $dt=1
M365 141 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=44670 $dt=1
M366 140 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=45530 $dt=1
M367 139 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=49210 $dt=1
M368 10 71 146 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=31910 $dt=1
M369 10 71 145 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=35590 $dt=1
M370 10 71 144 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=36450 $dt=1
M371 10 71 143 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40130 $dt=1
M372 10 71 142 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40990 $dt=1
M373 10 71 141 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=44670 $dt=1
M374 10 71 140 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=45530 $dt=1
M375 10 71 139 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=49210 $dt=1
M376 80 146 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=31860 $dt=1
M377 81 145 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=35400 $dt=1
M378 82 144 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=36400 $dt=1
M379 75 143 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=39940 $dt=1
M380 76 142 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=40940 $dt=1
M381 77 141 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=44480 $dt=1
M382 78 140 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=45480 $dt=1
M383 79 139 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=49020 $dt=1
.ends WallaceMultiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055847                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055847 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055847

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055819                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055819 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7655933055819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055820                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055820 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7655933055820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055821                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055821 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7655933055821

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055822                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055822 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7655933055822

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7655933055823                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7655933055823 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7655933055823

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055824                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055824 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.6986 scb=0.0347897 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7655933055824

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055825                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055825 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7655933055825

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055826                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055826 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7655933055826

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7655933055827                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7655933055827 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7655933055827

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAdder 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=10
X0 8 M2_M1_CDNS_765593305586 $T=2700 5110 0 90 $X=2570 $Y=5030
X1 9 M2_M1_CDNS_765593305586 $T=3060 2950 0 90 $X=2930 $Y=2870
X2 9 M2_M1_CDNS_765593305586 $T=3060 5520 0 90 $X=2930 $Y=5440
X3 5 M2_M1_CDNS_765593305586 $T=3450 7370 0 90 $X=3320 $Y=7290
X4 3 M2_M1_CDNS_765593305586 $T=3450 8190 0 90 $X=3320 $Y=8110
X5 5 M2_M1_CDNS_765593305586 $T=3460 3880 0 90 $X=3330 $Y=3800
X6 3 M2_M1_CDNS_765593305586 $T=4250 4700 0 90 $X=4120 $Y=4620
X7 10 M2_M1_CDNS_765593305586 $T=4700 5110 0 90 $X=4570 $Y=5030
X8 10 M2_M1_CDNS_765593305586 $T=4740 5820 0 90 $X=4610 $Y=5740
X9 8 M2_M1_CDNS_765593305586 $T=5140 5990 0 90 $X=5010 $Y=5910
X10 8 M2_M1_CDNS_765593305588 $T=5020 6720 0 90 $X=4890 $Y=6590
X11 10 M1_PO_CDNS_7655933055841 $T=1550 6040 0 90 $X=1430 $Y=5940
X12 5 M1_PO_CDNS_7655933055841 $T=3090 2650 0 90 $X=2970 $Y=2550
X13 5 M1_PO_CDNS_7655933055841 $T=3090 3820 0 90 $X=2970 $Y=3720
X14 5 M1_PO_CDNS_7655933055841 $T=3090 4360 0 90 $X=2970 $Y=4260
X15 6 M1_PO_CDNS_7655933055841 $T=3145 6870 0 90 $X=3025 $Y=6770
X16 9 M1_PO_CDNS_7655933055841 $T=3720 5020 0 90 $X=3600 $Y=4920
X17 8 M2_M1_CDNS_7655933055843 $T=2700 7470 0 90 $X=2450 $Y=7390
X18 6 M2_M1_CDNS_7655933055843 $T=3820 6180 0 90 $X=3570 $Y=6100
X19 3 M2_M1_CDNS_7655933055843 $T=4200 5220 0 90 $X=3950 $Y=5140
X20 3 M2_M1_CDNS_7655933055843 $T=4250 4170 0 90 $X=4000 $Y=4090
X21 10 M2_M1_CDNS_7655933055843 $T=4650 8090 0 90 $X=4400 $Y=8010
X22 8 M1_PO_CDNS_7655933055844 $T=2700 7470 0 90 $X=2450 $Y=7370
X23 6 M1_PO_CDNS_7655933055844 $T=3820 6180 0 90 $X=3570 $Y=6080
X24 3 M1_PO_CDNS_7655933055844 $T=4200 5220 0 90 $X=3950 $Y=5120
X25 3 M1_PO_CDNS_7655933055844 $T=4250 4170 0 90 $X=4000 $Y=4070
X26 10 M1_PO_CDNS_7655933055844 $T=4650 8090 0 90 $X=4400 $Y=7990
X27 8 M1_PO_CDNS_7655933055844 $T=5020 6720 0 90 $X=4770 $Y=6620
X28 9 3 8 1 nmos1v_CDNS_765593305588 $T=2220 5270 0 90 $X=1780 $Y=5030
X29 10 6 2 1 nmos1v_CDNS_765593305588 $T=2220 6290 1 270 $X=1780 $Y=5780
X30 3 10 4 1 nmos1v_CDNS_765593305588 $T=2220 7950 0 90 $X=1780 $Y=7710
X31 5 3 8 1 7 pmos1v_CDNS_7655933055812 $T=5670 4040 0 90 $X=5230 $Y=3620
X32 9 3 10 1 7 pmos1v_CDNS_7655933055812 $T=5670 5360 1 270 $X=5230 $Y=5030
X33 5 8 4 1 7 pmos1v_CDNS_7655933055812 $T=5670 7540 0 90 $X=5230 $Y=7120
X34 6 M2_M1_CDNS_7655933055847 $T=3820 2110 0 90 $X=3740 $Y=1860
X35 3 M2_M1_CDNS_7655933055847 $T=4260 2110 0 90 $X=4180 $Y=1860
X36 1 1 5 9 nmos1v_CDNS_7655933055819 $T=2220 3200 1 270 $X=1420 $Y=2690
X37 5 3 10 1 nmos1v_CDNS_7655933055820 $T=2220 4450 0 90 $X=1780 $Y=4210
X38 10 5 3 1 nmos1v_CDNS_7655933055821 $T=2220 4130 1 270 $X=1780 $Y=3620
X39 2 6 10 1 nmos1v_CDNS_7655933055821 $T=2220 6610 0 90 $X=1780 $Y=6250
X40 4 6 8 1 nmos1v_CDNS_7655933055821 $T=2220 7630 1 270 $X=1780 $Y=7120
X41 6 8 2 1 7 pmos1v_CDNS_7655933055822 $T=5670 6700 1 270 $X=5230 $Y=6250
X42 6 10 4 1 7 pmos1v_CDNS_7655933055822 $T=5670 8040 1 270 $X=5230 $Y=7590
X43 8 3 9 1 nmos1v_CDNS_7655933055823 $T=2220 4950 1 270 $X=1780 $Y=4500
X44 8 5 3 1 7 pmos1v_CDNS_7655933055824 $T=5670 4540 1 270 $X=5230 $Y=4090
X45 3 10 9 1 7 pmos1v_CDNS_7655933055825 $T=5670 4860 0 90 $X=5230 $Y=4500
X46 7 7 5 9 1 pmos1v_CDNS_7655933055826 $T=5670 3200 1 270 $X=5230 $Y=2690
X47 8 6 2 1 7 pmos1v_CDNS_7655933055827 $T=5670 6200 0 90 $X=5230 $Y=5780
M0 4 8 6 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=7540 $dt=0
M1 7 5 9 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5430 $Y=3110 $dt=1
M2 8 3 5 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5430 $Y=4040 $dt=1
M3 9 3 10 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5430 $Y=5270 $dt=1
M4 6 8 2 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=95.6709 scb=0.0347795 scc=0.0111862 $X=5430 $Y=6610 $dt=1
M5 4 8 5 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=99.6807 scb=0.0402027 scc=0.0112574 $X=5430 $Y=7540 $dt=1
.ends FAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7655933055848                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7655933055848 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7655933055848

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055849                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055849 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055849

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055850                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055850 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055850

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055851                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055851 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055851

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055852                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055852 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055852

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055853                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055853 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055853

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7655933055854                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7655933055854 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7655933055854

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X0 6 M2_M1_CDNS_765593305586 $T=690 3330 0 0 $X=610 $Y=3200
X1 1 M2_M1_CDNS_765593305586 $T=1190 1490 0 0 $X=1110 $Y=1360
X2 1 M2_M1_CDNS_765593305586 $T=2520 1490 0 0 $X=2440 $Y=1360
X3 6 M2_M1_CDNS_765593305586 $T=2550 3330 0 0 $X=2470 $Y=3200
X4 7 M1_PO_CDNS_7655933055841 $T=2470 2570 0 0 $X=2370 $Y=2450
X5 2 2 1 6 3 pmos1v_CDNS_765593305580 $T=420 3660 0 0 $X=0 $Y=3460
X6 1 2 5 4 3 pmos1v_CDNS_765593305580 $T=1350 3660 0 0 $X=930 $Y=3460
X7 6 2 7 4 3 pmos1v_CDNS_765593305580 $T=2370 3660 1 180 $X=1860 $Y=3460
X8 2 2 5 7 3 pmos1v_CDNS_765593305580 $T=3300 3660 1 180 $X=2790 $Y=3460
X9 3 3 1 6 nmos1v_CDNS_765593305581 $T=420 800 0 0 $X=0 $Y=240
X10 4 3 5 6 nmos1v_CDNS_765593305581 $T=1440 800 1 180 $X=930 $Y=240
X11 4 3 7 1 nmos1v_CDNS_765593305581 $T=2280 800 0 0 $X=1860 $Y=240
X12 3 3 5 7 nmos1v_CDNS_765593305581 $T=3300 800 1 180 $X=2790 $Y=240
X13 1 M2_M1_CDNS_7655933055843 $T=320 1490 0 0 $X=240 $Y=1240
X14 5 M2_M1_CDNS_7655933055843 $T=1540 2050 0 0 $X=1460 $Y=1800
X15 5 M2_M1_CDNS_7655933055843 $T=3400 2050 0 0 $X=3320 $Y=1800
X16 1 M1_PO_CDNS_7655933055844 $T=320 1490 0 0 $X=220 $Y=1240
X17 5 M1_PO_CDNS_7655933055844 $T=1540 2050 0 0 $X=1440 $Y=1800
X18 5 M1_PO_CDNS_7655933055844 $T=3400 2050 0 0 $X=3300 $Y=1800
X19 4 M5_M4_CDNS_7655933055850 $T=1850 2810 0 90 $X=1600 $Y=2590
X20 4 M4_M3_CDNS_7655933055851 $T=1850 2810 0 90 $X=1600 $Y=2590
X21 4 M3_M2_CDNS_7655933055852 $T=1850 2810 0 90 $X=1600 $Y=2590
X22 4 M2_M1_CDNS_7655933055853 $T=1850 2810 0 90 $X=1600 $Y=2590
X23 4 M6_M5_CDNS_7655933055854 $T=1850 2810 0 90 $X=1600 $Y=2590
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=420 $Y=800 $dt=0
M1 4 5 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1350 $Y=800 $dt=0
M2 1 7 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=2280 $Y=800 $dt=0
M3 3 5 7 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=3210 $Y=800 $dt=0
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7655933055855                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7655933055855 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7655933055855

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7655933055856                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7655933055856 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7655933055856

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7655933055857                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7655933055857 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7655933055857

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7655933055858                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7655933055858 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7655933055858

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7655933055859                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7655933055859 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7655933055859

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7655933055861                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7655933055861 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7655933055861

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7655933055862                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7655933055862 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7655933055862

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7655933055863                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7655933055863 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7655933055863

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7655933055864                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7655933055864 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7655933055864

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7655933055865                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7655933055865 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7655933055865

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7655933055866                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7655933055866 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7655933055866

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39
*.DEVICECLIMB
** N=39 EP=39 FDC=54
X0 2 M2_M1_CDNS_765593305580 $T=610 4030 0 0 $X=530 $Y=3780
X1 1 M2_M1_CDNS_765593305580 $T=930 5440 0 0 $X=850 $Y=5190
X2 3 M2_M1_CDNS_765593305580 $T=1860 4970 0 0 $X=1780 $Y=4720
X3 2 M2_M1_CDNS_765593305580 $T=2790 4030 0 0 $X=2710 $Y=3780
X4 7 M2_M1_CDNS_765593305580 $T=3110 3560 0 0 $X=3030 $Y=3310
X5 8 M2_M1_CDNS_765593305580 $T=4110 1490 0 0 $X=4030 $Y=1240
X6 6 M2_M1_CDNS_765593305580 $T=4650 5910 0 0 $X=4570 $Y=5660
X7 1 M2_M1_CDNS_765593305580 $T=5580 5440 0 0 $X=5500 $Y=5190
X8 3 M2_M1_CDNS_765593305580 $T=6510 4970 0 0 $X=6430 $Y=4720
X9 2 M2_M1_CDNS_765593305580 $T=7440 4030 0 0 $X=7360 $Y=3780
X10 7 M2_M1_CDNS_765593305580 $T=8370 3560 0 0 $X=8290 $Y=3310
X11 10 M2_M1_CDNS_765593305580 $T=8700 3090 0 0 $X=8620 $Y=2840
X12 11 M2_M1_CDNS_765593305580 $T=9690 1490 0 0 $X=9610 $Y=1240
X13 9 M2_M1_CDNS_765593305580 $T=10230 6380 0 0 $X=10150 $Y=6130
X14 6 M2_M1_CDNS_765593305580 $T=11160 5910 0 0 $X=11080 $Y=5660
X15 1 M2_M1_CDNS_765593305580 $T=12090 5440 0 0 $X=12010 $Y=5190
X16 3 M2_M1_CDNS_765593305580 $T=13020 4970 0 0 $X=12940 $Y=4720
X17 2 M2_M1_CDNS_765593305580 $T=13950 4030 0 0 $X=13870 $Y=3780
X18 7 M2_M1_CDNS_765593305580 $T=14880 3560 0 0 $X=14800 $Y=3310
X19 10 M2_M1_CDNS_765593305580 $T=15810 3090 0 0 $X=15730 $Y=2840
X20 13 M2_M1_CDNS_765593305580 $T=17130 1490 0 0 $X=17050 $Y=1240
X21 14 M2_M1_CDNS_765593305580 $T=17490 2630 0 0 $X=17410 $Y=2380
X22 12 M2_M1_CDNS_765593305580 $T=17670 6850 0 0 $X=17590 $Y=6600
X23 9 M2_M1_CDNS_765593305580 $T=18600 6380 0 0 $X=18520 $Y=6130
X24 6 M2_M1_CDNS_765593305580 $T=19530 5910 0 0 $X=19450 $Y=5660
X25 1 M2_M1_CDNS_765593305580 $T=20460 5440 0 0 $X=20380 $Y=5190
X26 3 M2_M1_CDNS_765593305580 $T=21390 4970 0 0 $X=21310 $Y=4720
X27 2 M2_M1_CDNS_765593305580 $T=22320 4030 0 0 $X=22240 $Y=3780
X28 7 M2_M1_CDNS_765593305580 $T=23250 3560 0 0 $X=23170 $Y=3310
X29 10 M2_M1_CDNS_765593305580 $T=24180 3090 0 0 $X=24100 $Y=2840
X30 14 M2_M1_CDNS_765593305580 $T=25110 2620 0 0 $X=25030 $Y=2370
X31 15 M2_M1_CDNS_765593305580 $T=26430 1490 0 0 $X=26350 $Y=1240
X32 7 M4_M3_CDNS_765593305581 $T=3110 3560 0 0 $X=3030 $Y=3310
X33 8 M4_M3_CDNS_765593305581 $T=4110 1490 0 0 $X=4030 $Y=1240
X34 11 M4_M3_CDNS_765593305581 $T=9690 1490 0 0 $X=9610 $Y=1240
X35 13 M4_M3_CDNS_765593305581 $T=17130 1490 0 0 $X=17050 $Y=1240
X36 14 M4_M3_CDNS_765593305581 $T=17490 2630 0 0 $X=17410 $Y=2380
X37 15 M4_M3_CDNS_765593305581 $T=26430 1490 0 0 $X=26350 $Y=1240
X38 2 M3_M2_CDNS_765593305582 $T=610 4030 0 0 $X=530 $Y=3780
X39 1 M3_M2_CDNS_765593305582 $T=930 5440 0 0 $X=850 $Y=5190
X40 2 M3_M2_CDNS_765593305582 $T=2790 4030 0 0 $X=2710 $Y=3780
X41 7 M3_M2_CDNS_765593305582 $T=3110 3560 0 0 $X=3030 $Y=3310
X42 8 M3_M2_CDNS_765593305582 $T=4110 1490 0 0 $X=4030 $Y=1240
X43 1 M3_M2_CDNS_765593305582 $T=5580 5440 0 0 $X=5500 $Y=5190
X44 2 M3_M2_CDNS_765593305582 $T=7440 4030 0 0 $X=7360 $Y=3780
X45 10 M3_M2_CDNS_765593305582 $T=8700 3090 0 0 $X=8620 $Y=2840
X46 11 M3_M2_CDNS_765593305582 $T=9690 1490 0 0 $X=9610 $Y=1240
X47 9 M3_M2_CDNS_765593305582 $T=10230 6380 0 0 $X=10150 $Y=6130
X48 1 M3_M2_CDNS_765593305582 $T=12090 5440 0 0 $X=12010 $Y=5190
X49 2 M3_M2_CDNS_765593305582 $T=13950 4030 0 0 $X=13870 $Y=3780
X50 10 M3_M2_CDNS_765593305582 $T=15810 3090 0 0 $X=15730 $Y=2840
X51 13 M3_M2_CDNS_765593305582 $T=17130 1490 0 0 $X=17050 $Y=1240
X52 14 M3_M2_CDNS_765593305582 $T=17490 2630 0 0 $X=17410 $Y=2380
X53 9 M3_M2_CDNS_765593305582 $T=18600 6380 0 0 $X=18520 $Y=6130
X54 1 M3_M2_CDNS_765593305582 $T=20460 5440 0 0 $X=20380 $Y=5190
X55 2 M3_M2_CDNS_765593305582 $T=22320 4030 0 0 $X=22240 $Y=3780
X56 10 M3_M2_CDNS_765593305582 $T=24180 3090 0 0 $X=24100 $Y=2840
X57 15 M3_M2_CDNS_765593305582 $T=26430 1490 0 0 $X=26350 $Y=1240
X58 3 M3_M2_CDNS_765593305585 $T=250 4970 0 90 $X=0 $Y=4890
X59 3 M3_M2_CDNS_765593305585 $T=1860 4970 0 0 $X=1780 $Y=4720
X60 6 M3_M2_CDNS_765593305585 $T=4650 5910 0 0 $X=4570 $Y=5660
X61 3 M3_M2_CDNS_765593305585 $T=6510 4970 0 0 $X=6430 $Y=4720
X62 7 M3_M2_CDNS_765593305585 $T=8370 3560 0 0 $X=8290 $Y=3310
X63 6 M3_M2_CDNS_765593305585 $T=11160 5910 0 0 $X=11080 $Y=5660
X64 3 M3_M2_CDNS_765593305585 $T=13020 4970 0 0 $X=12940 $Y=4720
X65 7 M3_M2_CDNS_765593305585 $T=14880 3560 0 0 $X=14800 $Y=3310
X66 12 M3_M2_CDNS_765593305585 $T=17670 6850 0 0 $X=17590 $Y=6600
X67 6 M3_M2_CDNS_765593305585 $T=19530 5910 0 0 $X=19450 $Y=5660
X68 3 M3_M2_CDNS_765593305585 $T=21390 4970 0 0 $X=21310 $Y=4720
X69 7 M3_M2_CDNS_765593305585 $T=23250 3560 0 0 $X=23170 $Y=3310
X70 14 M3_M2_CDNS_765593305585 $T=25110 2620 0 0 $X=25030 $Y=2370
X71 2 M5_M4_CDNS_7655933055822 $T=610 4030 0 0 $X=530 $Y=3780
X72 1 M5_M4_CDNS_7655933055822 $T=930 5440 0 0 $X=850 $Y=5190
X73 2 M5_M4_CDNS_7655933055822 $T=2790 4030 0 0 $X=2710 $Y=3780
X74 1 M5_M4_CDNS_7655933055822 $T=5580 5440 0 0 $X=5500 $Y=5190
X75 2 M5_M4_CDNS_7655933055822 $T=7440 4030 0 0 $X=7360 $Y=3780
X76 10 M5_M4_CDNS_7655933055822 $T=8700 3090 0 0 $X=8620 $Y=2840
X77 9 M5_M4_CDNS_7655933055822 $T=10230 6380 0 0 $X=10150 $Y=6130
X78 1 M5_M4_CDNS_7655933055822 $T=12090 5440 0 0 $X=12010 $Y=5190
X79 2 M5_M4_CDNS_7655933055822 $T=13950 4030 0 0 $X=13870 $Y=3780
X80 10 M5_M4_CDNS_7655933055822 $T=15810 3090 0 0 $X=15730 $Y=2840
X81 9 M5_M4_CDNS_7655933055822 $T=18600 6380 0 0 $X=18520 $Y=6130
X82 1 M5_M4_CDNS_7655933055822 $T=20460 5440 0 0 $X=20380 $Y=5190
X83 2 M5_M4_CDNS_7655933055822 $T=22320 4030 0 0 $X=22240 $Y=3780
X84 10 M5_M4_CDNS_7655933055822 $T=24180 3090 0 0 $X=24100 $Y=2840
X85 3 M2_M1_CDNS_7655933055829 $T=250 4970 0 90 $X=0 $Y=4890
X86 2 M4_M3_CDNS_7655933055836 $T=610 4030 0 0 $X=530 $Y=3780
X87 1 M4_M3_CDNS_7655933055836 $T=930 5440 0 0 $X=850 $Y=5190
X88 2 M4_M3_CDNS_7655933055836 $T=2790 4030 0 0 $X=2710 $Y=3780
X89 1 M4_M3_CDNS_7655933055836 $T=5580 5440 0 0 $X=5500 $Y=5190
X90 2 M4_M3_CDNS_7655933055836 $T=7440 4030 0 0 $X=7360 $Y=3780
X91 10 M4_M3_CDNS_7655933055836 $T=8700 3090 0 0 $X=8620 $Y=2840
X92 9 M4_M3_CDNS_7655933055836 $T=10230 6380 0 0 $X=10150 $Y=6130
X93 1 M4_M3_CDNS_7655933055836 $T=12090 5440 0 0 $X=12010 $Y=5190
X94 2 M4_M3_CDNS_7655933055836 $T=13950 4030 0 0 $X=13870 $Y=3780
X95 10 M4_M3_CDNS_7655933055836 $T=15810 3090 0 0 $X=15730 $Y=2840
X96 9 M4_M3_CDNS_7655933055836 $T=18600 6380 0 0 $X=18520 $Y=6130
X97 1 M4_M3_CDNS_7655933055836 $T=20460 5440 0 0 $X=20380 $Y=5190
X98 2 M4_M3_CDNS_7655933055836 $T=22320 4030 0 0 $X=22240 $Y=3780
X99 10 M4_M3_CDNS_7655933055836 $T=24180 3090 0 0 $X=24100 $Y=2840
X100 4 4 2 16 5 pmos1v_CDNS_765593305580 $T=2980 8370 1 180 $X=2470 $Y=8170
X101 4 4 17 8 5 pmos1v_CDNS_765593305580 $T=3820 8370 0 0 $X=3400 $Y=8170
X102 4 4 6 18 5 pmos1v_CDNS_765593305580 $T=4750 8370 0 0 $X=4330 $Y=8170
X103 19 4 3 18 5 pmos1v_CDNS_765593305580 $T=6700 8370 1 180 $X=6190 $Y=8170
X104 20 4 2 19 5 pmos1v_CDNS_765593305580 $T=7630 8370 1 180 $X=7120 $Y=8170
X105 4 4 7 20 5 pmos1v_CDNS_765593305580 $T=8560 8370 1 180 $X=8050 $Y=8170
X106 4 4 18 11 5 pmos1v_CDNS_765593305580 $T=9400 8370 0 0 $X=8980 $Y=8170
X107 4 4 9 21 5 pmos1v_CDNS_765593305580 $T=10330 8370 0 0 $X=9910 $Y=8170
X108 22 4 6 21 5 pmos1v_CDNS_765593305580 $T=11350 8370 1 180 $X=10840 $Y=8170
X109 23 4 1 21 5 pmos1v_CDNS_765593305580 $T=12280 8370 1 180 $X=11770 $Y=8170
X110 24 4 3 21 5 pmos1v_CDNS_765593305580 $T=13210 8370 1 180 $X=12700 $Y=8170
X111 23 4 2 24 5 pmos1v_CDNS_765593305580 $T=14140 8370 1 180 $X=13630 $Y=8170
X112 22 4 7 23 5 pmos1v_CDNS_765593305580 $T=15070 8370 1 180 $X=14560 $Y=8170
X113 4 4 10 22 5 pmos1v_CDNS_765593305580 $T=16000 8370 1 180 $X=15490 $Y=8170
X114 4 4 12 25 5 pmos1v_CDNS_765593305580 $T=17770 8370 0 0 $X=17350 $Y=8170
X115 26 4 6 25 5 pmos1v_CDNS_765593305580 $T=19720 8370 1 180 $X=19210 $Y=8170
X116 27 4 1 25 5 pmos1v_CDNS_765593305580 $T=20650 8370 1 180 $X=20140 $Y=8170
X117 27 4 2 28 5 pmos1v_CDNS_765593305580 $T=22510 8370 1 180 $X=22000 $Y=8170
X118 26 4 7 27 5 pmos1v_CDNS_765593305580 $T=23440 8370 1 180 $X=22930 $Y=8170
X119 4 4 14 29 5 pmos1v_CDNS_765593305580 $T=25300 8370 1 180 $X=24790 $Y=8170
X120 4 4 25 15 5 pmos1v_CDNS_765593305580 $T=26140 8370 0 0 $X=25720 $Y=8170
X121 5 5 1 30 nmos1v_CDNS_765593305581 $T=1030 800 0 0 $X=610 $Y=240
X122 30 5 3 17 nmos1v_CDNS_765593305581 $T=1960 800 0 0 $X=1540 $Y=240
X123 5 5 6 31 nmos1v_CDNS_765593305581 $T=4750 800 0 0 $X=4330 $Y=240
X124 31 5 2 18 nmos1v_CDNS_765593305581 $T=7540 800 0 0 $X=7120 $Y=240
X125 5 5 7 18 nmos1v_CDNS_765593305581 $T=8560 800 1 180 $X=8050 $Y=240
X126 5 5 18 11 nmos1v_CDNS_765593305581 $T=9400 800 0 0 $X=8980 $Y=240
X127 32 5 1 33 nmos1v_CDNS_765593305581 $T=12190 800 0 0 $X=11770 $Y=240
X128 33 5 3 21 nmos1v_CDNS_765593305581 $T=13120 800 0 0 $X=12700 $Y=240
X129 34 5 7 21 nmos1v_CDNS_765593305581 $T=14980 800 0 0 $X=14560 $Y=240
X130 5 5 10 21 nmos1v_CDNS_765593305581 $T=16000 800 1 180 $X=15490 $Y=240
X131 5 5 21 13 nmos1v_CDNS_765593305581 $T=16840 800 0 0 $X=16420 $Y=240
X132 35 5 9 36 nmos1v_CDNS_765593305581 $T=18700 800 0 0 $X=18280 $Y=240
X133 36 5 7 25 nmos1v_CDNS_765593305581 $T=23350 800 0 0 $X=22930 $Y=240
X134 5 5 25 15 nmos1v_CDNS_765593305581 $T=26140 800 0 0 $X=25720 $Y=240
X135 5 5 2 17 nmos1v_CDNS_7655933055819 $T=2980 1040 0 180 $X=2470 $Y=240
X136 5 5 17 8 nmos1v_CDNS_7655933055819 $T=3820 1040 1 0 $X=3400 $Y=240
X137 31 5 1 37 nmos1v_CDNS_7655933055819 $T=5680 1040 1 0 $X=5260 $Y=240
X138 37 5 3 18 nmos1v_CDNS_7655933055819 $T=6610 1040 1 0 $X=6190 $Y=240
X139 5 5 9 34 nmos1v_CDNS_7655933055819 $T=10330 1040 1 0 $X=9910 $Y=240
X140 34 5 6 32 nmos1v_CDNS_7655933055819 $T=11260 1040 1 0 $X=10840 $Y=240
X141 32 5 2 21 nmos1v_CDNS_7655933055819 $T=14050 1040 1 0 $X=13630 $Y=240
X142 5 5 12 35 nmos1v_CDNS_7655933055819 $T=17770 1040 1 0 $X=17350 $Y=240
X143 36 5 6 38 nmos1v_CDNS_7655933055819 $T=19630 1040 1 0 $X=19210 $Y=240
X144 38 5 1 39 nmos1v_CDNS_7655933055819 $T=20560 1040 1 0 $X=20140 $Y=240
X145 39 5 3 25 nmos1v_CDNS_7655933055819 $T=21490 1040 1 0 $X=21070 $Y=240
X146 38 5 2 25 nmos1v_CDNS_7655933055819 $T=22420 1040 1 0 $X=22000 $Y=240
X147 35 5 10 25 nmos1v_CDNS_7655933055819 $T=24280 1040 1 0 $X=23860 $Y=240
X148 5 5 14 25 nmos1v_CDNS_7655933055819 $T=25300 1040 0 180 $X=24790 $Y=240
X149 4 4 1 17 5 pmos1v_CDNS_7655933055826 $T=1030 8610 1 0 $X=610 $Y=8170
X150 16 4 3 17 5 pmos1v_CDNS_7655933055826 $T=2050 8610 0 180 $X=1540 $Y=8170
X151 20 4 1 18 5 pmos1v_CDNS_7655933055826 $T=5770 8610 0 180 $X=5260 $Y=8170
X152 4 4 21 13 5 pmos1v_CDNS_7655933055826 $T=16840 8610 1 0 $X=16420 $Y=8170
X153 29 4 9 25 5 pmos1v_CDNS_7655933055826 $T=18790 8610 0 180 $X=18280 $Y=8170
X154 28 4 3 25 5 pmos1v_CDNS_7655933055826 $T=21580 8610 0 180 $X=21070 $Y=8170
X155 29 4 10 26 5 pmos1v_CDNS_7655933055826 $T=24370 8610 0 180 $X=23860 $Y=8170
X156 17 M5_M4_CDNS_7655933055850 $T=3580 4500 0 0 $X=3360 $Y=4250
X157 18 M5_M4_CDNS_7655933055850 $T=9160 4500 0 0 $X=8940 $Y=4250
X158 21 M5_M4_CDNS_7655933055850 $T=16600 4500 0 0 $X=16380 $Y=4250
X159 25 M5_M4_CDNS_7655933055850 $T=25900 4500 0 0 $X=25680 $Y=4250
X160 17 M4_M3_CDNS_7655933055851 $T=3580 4500 0 0 $X=3360 $Y=4250
X161 18 M4_M3_CDNS_7655933055851 $T=9160 4500 0 0 $X=8940 $Y=4250
X162 21 M4_M3_CDNS_7655933055851 $T=16600 4500 0 0 $X=16380 $Y=4250
X163 25 M4_M3_CDNS_7655933055851 $T=25900 4500 0 0 $X=25680 $Y=4250
X164 17 M3_M2_CDNS_7655933055852 $T=3580 4500 0 0 $X=3360 $Y=4250
X165 18 M3_M2_CDNS_7655933055852 $T=9160 4500 0 0 $X=8940 $Y=4250
X166 21 M3_M2_CDNS_7655933055852 $T=16600 4500 0 0 $X=16380 $Y=4250
X167 25 M3_M2_CDNS_7655933055852 $T=25900 4500 0 0 $X=25680 $Y=4250
X168 17 M2_M1_CDNS_7655933055853 $T=3580 4500 0 0 $X=3360 $Y=4250
X169 18 M2_M1_CDNS_7655933055853 $T=9160 4500 0 0 $X=8940 $Y=4250
X170 21 M2_M1_CDNS_7655933055853 $T=16600 4500 0 0 $X=16380 $Y=4250
X171 25 M2_M1_CDNS_7655933055853 $T=25900 4500 0 0 $X=25680 $Y=4250
X172 1 M4_M3_CDNS_7655933055855 $T=80 5580 0 0 $X=0 $Y=5190
X173 17 M4_M3_CDNS_7655933055855 $T=1540 7840 0 0 $X=1460 $Y=7450
X174 6 M4_M3_CDNS_7655933055855 $T=2130 6050 0 0 $X=2050 $Y=5660
X175 17 M4_M3_CDNS_7655933055855 $T=2470 1570 0 0 $X=2390 $Y=1180
X176 18 M4_M3_CDNS_7655933055855 $T=5260 7840 0 0 $X=5180 $Y=7450
X177 18 M4_M3_CDNS_7655933055855 $T=6450 7840 0 0 $X=6370 $Y=7450
X178 18 M4_M3_CDNS_7655933055855 $T=6860 1570 0 0 $X=6780 $Y=1180
X179 9 M4_M3_CDNS_7655933055855 $T=7710 6520 0 0 $X=7630 $Y=6130
X180 18 M4_M3_CDNS_7655933055855 $T=8050 1570 0 0 $X=7970 $Y=1180
X181 21 M4_M3_CDNS_7655933055855 $T=10840 7840 0 0 $X=10760 $Y=7450
X182 21 M4_M3_CDNS_7655933055855 $T=12030 7840 0 0 $X=11950 $Y=7450
X183 21 M4_M3_CDNS_7655933055855 $T=12960 7840 0 0 $X=12880 $Y=7450
X184 21 M4_M3_CDNS_7655933055855 $T=13370 1570 0 0 $X=13290 $Y=1180
X185 21 M4_M3_CDNS_7655933055855 $T=14300 1570 0 0 $X=14220 $Y=1180
X186 21 M4_M3_CDNS_7655933055855 $T=15490 1570 0 0 $X=15410 $Y=1180
X187 12 M4_M3_CDNS_7655933055855 $T=16080 6990 0 0 $X=16000 $Y=6600
X188 25 M4_M3_CDNS_7655933055855 $T=18280 7840 0 0 $X=18200 $Y=7450
X189 25 M4_M3_CDNS_7655933055855 $T=19470 7840 0 0 $X=19390 $Y=7450
X190 25 M4_M3_CDNS_7655933055855 $T=20400 7840 0 0 $X=20320 $Y=7450
X191 25 M4_M3_CDNS_7655933055855 $T=21330 7840 0 0 $X=21250 $Y=7450
X192 25 M4_M3_CDNS_7655933055855 $T=21740 1570 0 0 $X=21660 $Y=1180
X193 25 M4_M3_CDNS_7655933055855 $T=22670 1570 0 0 $X=22590 $Y=1180
X194 25 M4_M3_CDNS_7655933055855 $T=23600 1570 0 0 $X=23520 $Y=1180
X195 25 M4_M3_CDNS_7655933055855 $T=24790 1570 0 0 $X=24710 $Y=1180
X196 17 M7_M6_CDNS_7655933055856 $T=1540 7840 0 0 $X=1460 $Y=7450
X197 17 M7_M6_CDNS_7655933055856 $T=2470 1570 0 0 $X=2390 $Y=1180
X198 18 M7_M6_CDNS_7655933055856 $T=5260 7840 0 0 $X=5180 $Y=7450
X199 18 M7_M6_CDNS_7655933055856 $T=6450 7840 0 0 $X=6370 $Y=7450
X200 18 M7_M6_CDNS_7655933055856 $T=6860 1570 0 0 $X=6780 $Y=1180
X201 18 M7_M6_CDNS_7655933055856 $T=8050 1570 0 0 $X=7970 $Y=1180
X202 21 M7_M6_CDNS_7655933055856 $T=10840 7840 0 0 $X=10760 $Y=7450
X203 21 M7_M6_CDNS_7655933055856 $T=12030 7840 0 0 $X=11950 $Y=7450
X204 21 M7_M6_CDNS_7655933055856 $T=12960 7840 0 0 $X=12880 $Y=7450
X205 21 M7_M6_CDNS_7655933055856 $T=13370 1570 0 0 $X=13290 $Y=1180
X206 21 M7_M6_CDNS_7655933055856 $T=14300 1570 0 0 $X=14220 $Y=1180
X207 21 M7_M6_CDNS_7655933055856 $T=15490 1570 0 0 $X=15410 $Y=1180
X208 25 M7_M6_CDNS_7655933055856 $T=18280 7840 0 0 $X=18200 $Y=7450
X209 25 M7_M6_CDNS_7655933055856 $T=19470 7840 0 0 $X=19390 $Y=7450
X210 25 M7_M6_CDNS_7655933055856 $T=20400 7840 0 0 $X=20320 $Y=7450
X211 25 M7_M6_CDNS_7655933055856 $T=21330 7840 0 0 $X=21250 $Y=7450
X212 25 M7_M6_CDNS_7655933055856 $T=21740 1570 0 0 $X=21660 $Y=1180
X213 25 M7_M6_CDNS_7655933055856 $T=22670 1570 0 0 $X=22590 $Y=1180
X214 25 M7_M6_CDNS_7655933055856 $T=23600 1570 0 0 $X=23520 $Y=1180
X215 25 M7_M6_CDNS_7655933055856 $T=24790 1570 0 0 $X=24710 $Y=1180
X216 17 M1_PO_CDNS_7655933055857 $T=3580 4500 0 0 $X=3340 $Y=4250
X217 18 M1_PO_CDNS_7655933055857 $T=9160 4500 0 0 $X=8920 $Y=4250
X218 21 M1_PO_CDNS_7655933055857 $T=16600 4500 0 0 $X=16360 $Y=4250
X219 17 M6_M5_CDNS_7655933055858 $T=3580 4500 0 0 $X=3360 $Y=4250
X220 18 M6_M5_CDNS_7655933055858 $T=9160 4500 0 0 $X=8940 $Y=4250
X221 21 M6_M5_CDNS_7655933055858 $T=16600 4500 0 0 $X=16380 $Y=4250
X222 25 M6_M5_CDNS_7655933055858 $T=25900 4500 0 0 $X=25680 $Y=4250
X223 1 M1_PO_CDNS_7655933055859 $T=930 5440 0 0 $X=830 $Y=5190
X224 3 M1_PO_CDNS_7655933055859 $T=1860 4970 0 0 $X=1760 $Y=4720
X225 2 M1_PO_CDNS_7655933055859 $T=2790 4030 0 0 $X=2690 $Y=3780
X226 6 M1_PO_CDNS_7655933055859 $T=4650 5910 0 0 $X=4550 $Y=5660
X227 1 M1_PO_CDNS_7655933055859 $T=5580 5440 0 0 $X=5480 $Y=5190
X228 3 M1_PO_CDNS_7655933055859 $T=6510 4970 0 0 $X=6410 $Y=4720
X229 2 M1_PO_CDNS_7655933055859 $T=7440 4030 0 0 $X=7340 $Y=3780
X230 7 M1_PO_CDNS_7655933055859 $T=8370 3560 0 0 $X=8270 $Y=3310
X231 9 M1_PO_CDNS_7655933055859 $T=10230 6380 0 0 $X=10130 $Y=6130
X232 6 M1_PO_CDNS_7655933055859 $T=11160 5910 0 0 $X=11060 $Y=5660
X233 1 M1_PO_CDNS_7655933055859 $T=12090 5440 0 0 $X=11990 $Y=5190
X234 3 M1_PO_CDNS_7655933055859 $T=13020 4970 0 0 $X=12920 $Y=4720
X235 2 M1_PO_CDNS_7655933055859 $T=13950 4030 0 0 $X=13850 $Y=3780
X236 7 M1_PO_CDNS_7655933055859 $T=14880 3560 0 0 $X=14780 $Y=3310
X237 10 M1_PO_CDNS_7655933055859 $T=15810 3090 0 0 $X=15710 $Y=2840
X238 12 M1_PO_CDNS_7655933055859 $T=17670 6850 0 0 $X=17570 $Y=6600
X239 9 M1_PO_CDNS_7655933055859 $T=18600 6380 0 0 $X=18500 $Y=6130
X240 6 M1_PO_CDNS_7655933055859 $T=19530 5910 0 0 $X=19430 $Y=5660
X241 1 M1_PO_CDNS_7655933055859 $T=20460 5440 0 0 $X=20360 $Y=5190
X242 3 M1_PO_CDNS_7655933055859 $T=21390 4970 0 0 $X=21290 $Y=4720
X243 2 M1_PO_CDNS_7655933055859 $T=22320 4030 0 0 $X=22220 $Y=3780
X244 7 M1_PO_CDNS_7655933055859 $T=23250 3560 0 0 $X=23150 $Y=3310
X245 10 M1_PO_CDNS_7655933055859 $T=24180 3090 0 0 $X=24080 $Y=2840
X246 14 M1_PO_CDNS_7655933055859 $T=25110 2620 0 0 $X=25010 $Y=2370
X247 1 M2_M1_CDNS_7655933055861 $T=80 5580 0 0 $X=0 $Y=5190
X248 17 M2_M1_CDNS_7655933055861 $T=1540 7840 0 0 $X=1460 $Y=7450
X249 6 M2_M1_CDNS_7655933055861 $T=2130 6050 0 0 $X=2050 $Y=5660
X250 17 M2_M1_CDNS_7655933055861 $T=2470 1570 0 0 $X=2390 $Y=1180
X251 18 M2_M1_CDNS_7655933055861 $T=5260 7840 0 0 $X=5180 $Y=7450
X252 18 M2_M1_CDNS_7655933055861 $T=6450 7840 0 0 $X=6370 $Y=7450
X253 18 M2_M1_CDNS_7655933055861 $T=6860 1570 0 0 $X=6780 $Y=1180
X254 9 M2_M1_CDNS_7655933055861 $T=7710 6520 0 0 $X=7630 $Y=6130
X255 18 M2_M1_CDNS_7655933055861 $T=8050 1570 0 0 $X=7970 $Y=1180
X256 21 M2_M1_CDNS_7655933055861 $T=10840 7840 0 0 $X=10760 $Y=7450
X257 21 M2_M1_CDNS_7655933055861 $T=12030 7840 0 0 $X=11950 $Y=7450
X258 21 M2_M1_CDNS_7655933055861 $T=12960 7840 0 0 $X=12880 $Y=7450
X259 21 M2_M1_CDNS_7655933055861 $T=13370 1570 0 0 $X=13290 $Y=1180
X260 21 M2_M1_CDNS_7655933055861 $T=14300 1570 0 0 $X=14220 $Y=1180
X261 21 M2_M1_CDNS_7655933055861 $T=15490 1570 0 0 $X=15410 $Y=1180
X262 12 M2_M1_CDNS_7655933055861 $T=16080 6990 0 0 $X=16000 $Y=6600
X263 25 M2_M1_CDNS_7655933055861 $T=18280 7840 0 0 $X=18200 $Y=7450
X264 25 M2_M1_CDNS_7655933055861 $T=19470 7840 0 0 $X=19390 $Y=7450
X265 25 M2_M1_CDNS_7655933055861 $T=20400 7840 0 0 $X=20320 $Y=7450
X266 25 M2_M1_CDNS_7655933055861 $T=21330 7840 0 0 $X=21250 $Y=7450
X267 25 M2_M1_CDNS_7655933055861 $T=21740 1570 0 0 $X=21660 $Y=1180
X268 25 M2_M1_CDNS_7655933055861 $T=22670 1570 0 0 $X=22590 $Y=1180
X269 25 M2_M1_CDNS_7655933055861 $T=23600 1570 0 0 $X=23520 $Y=1180
X270 25 M2_M1_CDNS_7655933055861 $T=24790 1570 0 0 $X=24710 $Y=1180
X271 17 M7_M6_CDNS_7655933055862 $T=3580 4500 0 0 $X=3360 $Y=4250
X272 18 M7_M6_CDNS_7655933055862 $T=9160 4500 0 0 $X=8940 $Y=4250
X273 21 M7_M6_CDNS_7655933055862 $T=16600 4500 0 0 $X=16380 $Y=4250
X274 25 M7_M6_CDNS_7655933055862 $T=25900 4500 0 0 $X=25680 $Y=4250
X275 17 M6_M5_CDNS_7655933055863 $T=1540 7840 0 0 $X=1460 $Y=7450
X276 17 M6_M5_CDNS_7655933055863 $T=2470 1570 0 0 $X=2390 $Y=1180
X277 18 M6_M5_CDNS_7655933055863 $T=5260 7840 0 0 $X=5180 $Y=7450
X278 18 M6_M5_CDNS_7655933055863 $T=6450 7840 0 0 $X=6370 $Y=7450
X279 18 M6_M5_CDNS_7655933055863 $T=6860 1570 0 0 $X=6780 $Y=1180
X280 18 M6_M5_CDNS_7655933055863 $T=8050 1570 0 0 $X=7970 $Y=1180
X281 21 M6_M5_CDNS_7655933055863 $T=10840 7840 0 0 $X=10760 $Y=7450
X282 21 M6_M5_CDNS_7655933055863 $T=12030 7840 0 0 $X=11950 $Y=7450
X283 21 M6_M5_CDNS_7655933055863 $T=12960 7840 0 0 $X=12880 $Y=7450
X284 21 M6_M5_CDNS_7655933055863 $T=13370 1570 0 0 $X=13290 $Y=1180
X285 21 M6_M5_CDNS_7655933055863 $T=14300 1570 0 0 $X=14220 $Y=1180
X286 21 M6_M5_CDNS_7655933055863 $T=15490 1570 0 0 $X=15410 $Y=1180
X287 25 M6_M5_CDNS_7655933055863 $T=18280 7840 0 0 $X=18200 $Y=7450
X288 25 M6_M5_CDNS_7655933055863 $T=19470 7840 0 0 $X=19390 $Y=7450
X289 25 M6_M5_CDNS_7655933055863 $T=20400 7840 0 0 $X=20320 $Y=7450
X290 25 M6_M5_CDNS_7655933055863 $T=21330 7840 0 0 $X=21250 $Y=7450
X291 25 M6_M5_CDNS_7655933055863 $T=21740 1570 0 0 $X=21660 $Y=1180
X292 25 M6_M5_CDNS_7655933055863 $T=22670 1570 0 0 $X=22590 $Y=1180
X293 25 M6_M5_CDNS_7655933055863 $T=23600 1570 0 0 $X=23520 $Y=1180
X294 25 M6_M5_CDNS_7655933055863 $T=24790 1570 0 0 $X=24710 $Y=1180
X295 1 M6_M5_CDNS_7655933055864 $T=80 5580 0 0 $X=0 $Y=5190
X296 6 M6_M5_CDNS_7655933055864 $T=2130 6050 0 0 $X=2050 $Y=5660
X297 9 M6_M5_CDNS_7655933055864 $T=7710 6520 0 0 $X=7630 $Y=6130
X298 12 M6_M5_CDNS_7655933055864 $T=16080 6990 0 0 $X=16000 $Y=6600
X299 1 M3_M2_CDNS_7655933055865 $T=80 5580 0 0 $X=0 $Y=5190
X300 17 M3_M2_CDNS_7655933055865 $T=1540 7840 0 0 $X=1460 $Y=7450
X301 6 M3_M2_CDNS_7655933055865 $T=2130 6050 0 0 $X=2050 $Y=5660
X302 17 M3_M2_CDNS_7655933055865 $T=2470 1570 0 0 $X=2390 $Y=1180
X303 18 M3_M2_CDNS_7655933055865 $T=5260 7840 0 0 $X=5180 $Y=7450
X304 18 M3_M2_CDNS_7655933055865 $T=6450 7840 0 0 $X=6370 $Y=7450
X305 18 M3_M2_CDNS_7655933055865 $T=6860 1570 0 0 $X=6780 $Y=1180
X306 9 M3_M2_CDNS_7655933055865 $T=7710 6520 0 0 $X=7630 $Y=6130
X307 18 M3_M2_CDNS_7655933055865 $T=8050 1570 0 0 $X=7970 $Y=1180
X308 21 M3_M2_CDNS_7655933055865 $T=10840 7840 0 0 $X=10760 $Y=7450
X309 21 M3_M2_CDNS_7655933055865 $T=12030 7840 0 0 $X=11950 $Y=7450
X310 21 M3_M2_CDNS_7655933055865 $T=12960 7840 0 0 $X=12880 $Y=7450
X311 21 M3_M2_CDNS_7655933055865 $T=13370 1570 0 0 $X=13290 $Y=1180
X312 21 M3_M2_CDNS_7655933055865 $T=14300 1570 0 0 $X=14220 $Y=1180
X313 21 M3_M2_CDNS_7655933055865 $T=15490 1570 0 0 $X=15410 $Y=1180
X314 12 M3_M2_CDNS_7655933055865 $T=16080 6990 0 0 $X=16000 $Y=6600
X315 25 M3_M2_CDNS_7655933055865 $T=18280 7840 0 0 $X=18200 $Y=7450
X316 25 M3_M2_CDNS_7655933055865 $T=19470 7840 0 0 $X=19390 $Y=7450
X317 25 M3_M2_CDNS_7655933055865 $T=20400 7840 0 0 $X=20320 $Y=7450
X318 25 M3_M2_CDNS_7655933055865 $T=21330 7840 0 0 $X=21250 $Y=7450
X319 25 M3_M2_CDNS_7655933055865 $T=21740 1570 0 0 $X=21660 $Y=1180
X320 25 M3_M2_CDNS_7655933055865 $T=22670 1570 0 0 $X=22590 $Y=1180
X321 25 M3_M2_CDNS_7655933055865 $T=23600 1570 0 0 $X=23520 $Y=1180
X322 25 M3_M2_CDNS_7655933055865 $T=24790 1570 0 0 $X=24710 $Y=1180
X323 1 M5_M4_CDNS_7655933055866 $T=80 5580 0 0 $X=0 $Y=5190
X324 17 M5_M4_CDNS_7655933055866 $T=1540 7840 0 0 $X=1460 $Y=7450
X325 6 M5_M4_CDNS_7655933055866 $T=2130 6050 0 0 $X=2050 $Y=5660
X326 17 M5_M4_CDNS_7655933055866 $T=2470 1570 0 0 $X=2390 $Y=1180
X327 18 M5_M4_CDNS_7655933055866 $T=5260 7840 0 0 $X=5180 $Y=7450
X328 18 M5_M4_CDNS_7655933055866 $T=6450 7840 0 0 $X=6370 $Y=7450
X329 18 M5_M4_CDNS_7655933055866 $T=6860 1570 0 0 $X=6780 $Y=1180
X330 9 M5_M4_CDNS_7655933055866 $T=7710 6520 0 0 $X=7630 $Y=6130
X331 18 M5_M4_CDNS_7655933055866 $T=8050 1570 0 0 $X=7970 $Y=1180
X332 21 M5_M4_CDNS_7655933055866 $T=10840 7840 0 0 $X=10760 $Y=7450
X333 21 M5_M4_CDNS_7655933055866 $T=12030 7840 0 0 $X=11950 $Y=7450
X334 21 M5_M4_CDNS_7655933055866 $T=12960 7840 0 0 $X=12880 $Y=7450
X335 21 M5_M4_CDNS_7655933055866 $T=13370 1570 0 0 $X=13290 $Y=1180
X336 21 M5_M4_CDNS_7655933055866 $T=14300 1570 0 0 $X=14220 $Y=1180
X337 21 M5_M4_CDNS_7655933055866 $T=15490 1570 0 0 $X=15410 $Y=1180
X338 12 M5_M4_CDNS_7655933055866 $T=16080 6990 0 0 $X=16000 $Y=6600
X339 25 M5_M4_CDNS_7655933055866 $T=18280 7840 0 0 $X=18200 $Y=7450
X340 25 M5_M4_CDNS_7655933055866 $T=19470 7840 0 0 $X=19390 $Y=7450
X341 25 M5_M4_CDNS_7655933055866 $T=20400 7840 0 0 $X=20320 $Y=7450
X342 25 M5_M4_CDNS_7655933055866 $T=21330 7840 0 0 $X=21250 $Y=7450
X343 25 M5_M4_CDNS_7655933055866 $T=21740 1570 0 0 $X=21660 $Y=1180
X344 25 M5_M4_CDNS_7655933055866 $T=22670 1570 0 0 $X=22590 $Y=1180
X345 25 M5_M4_CDNS_7655933055866 $T=23600 1570 0 0 $X=23520 $Y=1180
X346 25 M5_M4_CDNS_7655933055866 $T=24790 1570 0 0 $X=24710 $Y=1180
M0 30 1 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1030 $Y=800 $dt=0
M1 17 3 30 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1960 $Y=800 $dt=0
M2 31 6 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=4750 $Y=800 $dt=0
M3 18 2 31 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=7540 $Y=800 $dt=0
M4 5 7 18 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=8470 $Y=800 $dt=0
M5 11 18 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=9400 $Y=800 $dt=0
M6 33 1 32 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12190 $Y=800 $dt=0
M7 21 3 33 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=13120 $Y=800 $dt=0
M8 21 7 34 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=14980 $Y=800 $dt=0
M9 5 10 21 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=15910 $Y=800 $dt=0
M10 13 21 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=16840 $Y=800 $dt=0
M11 36 9 35 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=18700 $Y=800 $dt=0
M12 25 7 36 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=23350 $Y=800 $dt=0
M13 15 25 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=26140 $Y=800 $dt=0
M14 17 1 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=1030 $Y=8370 $dt=1
M15 16 3 17 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=1960 $Y=8370 $dt=1
M16 4 2 16 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M17 8 17 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M18 18 6 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M19 20 1 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=5680 $Y=8370 $dt=1
M20 19 3 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M21 20 2 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M22 4 7 20 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M23 11 18 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M24 21 9 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M25 22 6 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M26 23 1 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M27 24 3 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M28 23 2 24 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M29 22 7 23 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M30 4 10 22 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M31 13 21 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=16840 $Y=8370 $dt=1
M32 25 12 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M33 29 9 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=18700 $Y=8370 $dt=1
M34 26 6 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M35 27 1 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M36 28 3 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=21490 $Y=8370 $dt=1
M37 27 2 28 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M38 26 7 27 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
M39 29 10 26 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=24280 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceFinalAdder                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceFinalAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58
** N=164 EP=58 FDC=320
X0 33 M4_M3_CDNS_765593305581 $T=560 3210 0 0 $X=480 $Y=2960
X1 34 M4_M3_CDNS_765593305581 $T=9840 3210 0 0 $X=9760 $Y=2960
X2 35 M4_M3_CDNS_765593305581 $T=17280 3210 0 0 $X=17200 $Y=2960
X3 36 M4_M3_CDNS_765593305581 $T=22860 3210 0 0 $X=22780 $Y=2960
X4 37 M4_M3_CDNS_765593305581 $T=27230 3210 0 0 $X=27150 $Y=2960
X5 38 M4_M3_CDNS_765593305581 $T=36530 3210 0 0 $X=36450 $Y=2960
X6 39 M4_M3_CDNS_765593305581 $T=43970 3210 0 0 $X=43890 $Y=2960
X7 40 M4_M3_CDNS_765593305581 $T=49550 3210 0 0 $X=49470 $Y=2960
X8 41 M3_M2_CDNS_765593305582 $T=150 2650 0 0 $X=70 $Y=2400
X9 42 M3_M2_CDNS_765593305582 $T=5940 2650 0 0 $X=5860 $Y=2400
X10 43 M3_M2_CDNS_765593305582 $T=16170 2650 0 0 $X=16090 $Y=2400
X11 44 M3_M2_CDNS_765593305582 $T=21750 2650 0 0 $X=21670 $Y=2400
X12 45 M3_M2_CDNS_765593305582 $T=26890 2650 0 0 $X=26810 $Y=2400
X13 46 M3_M2_CDNS_765593305582 $T=32670 2650 0 0 $X=32590 $Y=2400
X14 47 M3_M2_CDNS_765593305582 $T=40090 2650 0 0 $X=40010 $Y=2400
X15 48 M3_M2_CDNS_765593305582 $T=48440 2650 0 0 $X=48360 $Y=2400
X16 49 M3_M2_CDNS_765593305582 $T=53580 2650 0 0 $X=53500 $Y=2400
X17 1 M2_M1_CDNS_765593305586 $T=4820 20240 0 0 $X=4740 $Y=20110
X18 9 M2_M1_CDNS_765593305586 $T=13610 20240 0 0 $X=13530 $Y=20110
X19 12 M2_M1_CDNS_765593305586 $T=19200 20240 0 0 $X=19120 $Y=20110
X20 17 M2_M1_CDNS_765593305586 $T=31060 20240 0 0 $X=30980 $Y=20110
X21 18 M2_M1_CDNS_765593305586 $T=31510 20240 0 0 $X=31430 $Y=20110
X22 21 M2_M1_CDNS_765593305586 $T=40300 20240 0 0 $X=40220 $Y=20110
X23 24 M2_M1_CDNS_765593305586 $T=45890 20240 0 0 $X=45810 $Y=20110
X24 30 M2_M1_CDNS_765593305586 $T=57710 20240 0 0 $X=57630 $Y=20110
X25 41 M4_M3_CDNS_7655933055836 $T=150 2650 0 0 $X=70 $Y=2400
X26 42 M4_M3_CDNS_7655933055836 $T=5940 2650 0 0 $X=5860 $Y=2400
X27 43 M4_M3_CDNS_7655933055836 $T=16170 2650 0 0 $X=16090 $Y=2400
X28 44 M4_M3_CDNS_7655933055836 $T=21750 2650 0 0 $X=21670 $Y=2400
X29 45 M4_M3_CDNS_7655933055836 $T=26890 2650 0 0 $X=26810 $Y=2400
X30 46 M4_M3_CDNS_7655933055836 $T=32670 2650 0 0 $X=32590 $Y=2400
X31 47 M4_M3_CDNS_7655933055836 $T=40090 2650 0 0 $X=40010 $Y=2400
X32 48 M4_M3_CDNS_7655933055836 $T=48440 2650 0 0 $X=48360 $Y=2400
X33 49 M4_M3_CDNS_7655933055836 $T=53580 2650 0 0 $X=53500 $Y=2400
X34 33 M3_M2_CDNS_7655933055838 $T=560 3210 0 0 $X=480 $Y=2960
X35 34 M3_M2_CDNS_7655933055838 $T=9840 3210 0 0 $X=9760 $Y=2960
X36 35 M3_M2_CDNS_7655933055838 $T=17280 3210 0 0 $X=17200 $Y=2960
X37 36 M3_M2_CDNS_7655933055838 $T=22860 3210 0 0 $X=22780 $Y=2960
X38 37 M3_M2_CDNS_7655933055838 $T=27230 3210 0 0 $X=27150 $Y=2960
X39 38 M3_M2_CDNS_7655933055838 $T=36530 3210 0 0 $X=36450 $Y=2960
X40 39 M3_M2_CDNS_7655933055838 $T=43970 3210 0 0 $X=43890 $Y=2960
X41 40 M3_M2_CDNS_7655933055838 $T=49550 3210 0 0 $X=49470 $Y=2960
X42 29 5 50 31 32 6 94 93 141 163
+ 164 142 HAdder $T=62720 6180 1 90 $X=53760 $Y=6980
X43 7 1 6 5 51 66 109 AND $T=3670 21910 0 0 $X=4740 $Y=18810
X44 10 9 6 5 52 70 112 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X45 13 12 6 5 53 73 115 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X46 15 17 6 5 54 80 128 AND $T=32210 21910 1 180 $X=26960 $Y=18810
X47 19 18 6 5 55 82 130 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X48 22 21 6 5 56 86 134 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X49 25 24 6 5 57 89 137 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X50 28 30 6 5 58 92 140 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X51 41 M6_M5_CDNS_7655933055848 $T=150 2650 0 0 $X=70 $Y=2400
X52 42 M6_M5_CDNS_7655933055848 $T=5940 2650 0 0 $X=5860 $Y=2400
X53 43 M6_M5_CDNS_7655933055848 $T=16170 2650 0 0 $X=16090 $Y=2400
X54 44 M6_M5_CDNS_7655933055848 $T=21750 2650 0 0 $X=21670 $Y=2400
X55 45 M6_M5_CDNS_7655933055848 $T=26890 2650 0 0 $X=26810 $Y=2400
X56 46 M6_M5_CDNS_7655933055848 $T=32670 2650 0 0 $X=32590 $Y=2400
X57 47 M6_M5_CDNS_7655933055848 $T=40090 2650 0 0 $X=40010 $Y=2400
X58 48 M6_M5_CDNS_7655933055848 $T=48440 2650 0 0 $X=48360 $Y=2400
X59 49 M6_M5_CDNS_7655933055848 $T=53580 2650 0 0 $X=53500 $Y=2400
X60 41 M5_M4_CDNS_7655933055849 $T=150 2650 0 0 $X=70 $Y=2400
X61 42 M5_M4_CDNS_7655933055849 $T=5940 2650 0 0 $X=5860 $Y=2400
X62 43 M5_M4_CDNS_7655933055849 $T=16170 2650 0 0 $X=16090 $Y=2400
X63 44 M5_M4_CDNS_7655933055849 $T=21750 2650 0 0 $X=21670 $Y=2400
X64 45 M5_M4_CDNS_7655933055849 $T=26890 2650 0 0 $X=26810 $Y=2400
X65 46 M5_M4_CDNS_7655933055849 $T=32670 2650 0 0 $X=32590 $Y=2400
X66 47 M5_M4_CDNS_7655933055849 $T=40090 2650 0 0 $X=40010 $Y=2400
X67 48 M5_M4_CDNS_7655933055849 $T=48440 2650 0 0 $X=48360 $Y=2400
X68 49 M5_M4_CDNS_7655933055849 $T=53580 2650 0 0 $X=53500 $Y=2400
X69 51 M5_M4_CDNS_7655933055850 $T=9340 19910 0 0 $X=9120 $Y=19660
X70 52 M5_M4_CDNS_7655933055850 $T=18130 19910 0 0 $X=17910 $Y=19660
X71 53 M5_M4_CDNS_7655933055850 $T=23720 19910 0 0 $X=23500 $Y=19660
X72 54 M5_M4_CDNS_7655933055850 $T=26500 19910 0 0 $X=26280 $Y=19660
X73 55 M5_M4_CDNS_7655933055850 $T=36030 19910 0 0 $X=35810 $Y=19660
X74 56 M5_M4_CDNS_7655933055850 $T=44820 19910 0 0 $X=44600 $Y=19660
X75 57 M5_M4_CDNS_7655933055850 $T=50410 19910 0 0 $X=50190 $Y=19660
X76 58 M5_M4_CDNS_7655933055850 $T=53190 19910 0 0 $X=52970 $Y=19660
X77 51 M4_M3_CDNS_7655933055851 $T=9340 19910 0 0 $X=9120 $Y=19660
X78 52 M4_M3_CDNS_7655933055851 $T=18130 19910 0 0 $X=17910 $Y=19660
X79 53 M4_M3_CDNS_7655933055851 $T=23720 19910 0 0 $X=23500 $Y=19660
X80 54 M4_M3_CDNS_7655933055851 $T=26500 19910 0 0 $X=26280 $Y=19660
X81 55 M4_M3_CDNS_7655933055851 $T=36030 19910 0 0 $X=35810 $Y=19660
X82 56 M4_M3_CDNS_7655933055851 $T=44820 19910 0 0 $X=44600 $Y=19660
X83 57 M4_M3_CDNS_7655933055851 $T=50410 19910 0 0 $X=50190 $Y=19660
X84 58 M4_M3_CDNS_7655933055851 $T=53190 19910 0 0 $X=52970 $Y=19660
X85 51 M3_M2_CDNS_7655933055852 $T=9340 19910 0 0 $X=9120 $Y=19660
X86 52 M3_M2_CDNS_7655933055852 $T=18130 19910 0 0 $X=17910 $Y=19660
X87 53 M3_M2_CDNS_7655933055852 $T=23720 19910 0 0 $X=23500 $Y=19660
X88 54 M3_M2_CDNS_7655933055852 $T=26500 19910 0 0 $X=26280 $Y=19660
X89 55 M3_M2_CDNS_7655933055852 $T=36030 19910 0 0 $X=35810 $Y=19660
X90 56 M3_M2_CDNS_7655933055852 $T=44820 19910 0 0 $X=44600 $Y=19660
X91 57 M3_M2_CDNS_7655933055852 $T=50410 19910 0 0 $X=50190 $Y=19660
X92 58 M3_M2_CDNS_7655933055852 $T=53190 19910 0 0 $X=52970 $Y=19660
X93 51 M2_M1_CDNS_7655933055853 $T=9340 19910 0 0 $X=9120 $Y=19660
X94 52 M2_M1_CDNS_7655933055853 $T=18130 19910 0 0 $X=17910 $Y=19660
X95 53 M2_M1_CDNS_7655933055853 $T=23720 19910 0 0 $X=23500 $Y=19660
X96 54 M2_M1_CDNS_7655933055853 $T=26500 19910 0 0 $X=26280 $Y=19660
X97 55 M2_M1_CDNS_7655933055853 $T=36030 19910 0 0 $X=35810 $Y=19660
X98 56 M2_M1_CDNS_7655933055853 $T=44820 19910 0 0 $X=44600 $Y=19660
X99 57 M2_M1_CDNS_7655933055853 $T=50410 19910 0 0 $X=50190 $Y=19660
X100 58 M2_M1_CDNS_7655933055853 $T=53190 19910 0 0 $X=52970 $Y=19660
X101 51 M6_M5_CDNS_7655933055854 $T=9340 19910 0 0 $X=9120 $Y=19660
X102 52 M6_M5_CDNS_7655933055854 $T=18130 19910 0 0 $X=17910 $Y=19660
X103 53 M6_M5_CDNS_7655933055854 $T=23720 19910 0 0 $X=23500 $Y=19660
X104 54 M6_M5_CDNS_7655933055854 $T=26500 19910 0 0 $X=26280 $Y=19660
X105 55 M6_M5_CDNS_7655933055854 $T=36030 19910 0 0 $X=35810 $Y=19660
X106 56 M6_M5_CDNS_7655933055854 $T=44820 19910 0 0 $X=44600 $Y=19660
X107 57 M6_M5_CDNS_7655933055854 $T=50410 19910 0 0 $X=50190 $Y=19660
X108 58 M6_M5_CDNS_7655933055854 $T=53190 19910 0 0 $X=52970 $Y=19660
X109 3 6 5 41 2 106 64 XOR $T=530 18810 1 0 $X=530 $Y=14110
X110 33 6 5 4 41 105 63 XOR $T=640 4700 1 0 $X=640 $Y=0
X111 1 6 5 42 7 108 65 XOR $T=4740 18810 1 0 $X=4740 $Y=14110
X112 34 6 5 8 42 107 67 XOR $T=9740 4700 0 180 $X=6020 $Y=0
X113 35 6 5 11 43 111 69 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X114 9 6 5 43 10 110 68 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X115 36 6 5 14 44 114 72 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X116 12 6 5 44 13 113 71 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X117 37 6 5 16 45 116 74 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X118 17 6 5 45 15 127 79 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X119 18 6 5 46 19 129 81 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X120 38 6 5 20 46 131 83 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X121 39 6 5 23 47 133 85 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X122 21 6 5 47 22 132 84 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X123 40 6 5 27 48 136 88 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X124 24 6 5 48 25 135 87 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X125 50 6 5 26 49 138 90 XOR $T=49650 4700 1 0 $X=49650 $Y=0
X126 30 6 5 49 28 139 91 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X127 45 54 37 6 5 44 53 36 43 52
+ 35 42 34 51 33 143 59 60 145 144
+ 61 146 147 148 62 150 151 152 149 95
+ 96 99 100 98 101 102 97 103 104 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X128 49 58 50 6 5 48 57 40 47 56
+ 39 46 38 55 37 153 75 76 155 154
+ 77 156 157 158 78 160 161 162 159 117
+ 118 121 122 120 123 124 119 125 126 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
M0 109 1 66 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5600 $Y=19150 $dt=0
M1 5 7 109 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5810 $Y=19150 $dt=0
M2 51 66 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=8230 $Y=19140 $dt=0
M3 112 9 70 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=19150 $dt=0
M4 5 10 112 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=19150 $dt=0
M5 52 70 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=19140 $dt=0
M6 115 12 73 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=19150 $dt=0
M7 5 13 115 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=19150 $dt=0
M8 53 73 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=19140 $dt=0
M9 5 80 54 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27560 $Y=19140 $dt=0
M10 128 15 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29980 $Y=19150 $dt=0
M11 80 17 128 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30190 $Y=19150 $dt=0
M12 130 18 82 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=19150 $dt=0
M13 5 19 130 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=19150 $dt=0
M14 55 82 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=19140 $dt=0
M15 134 21 86 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=19150 $dt=0
M16 5 22 134 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=19150 $dt=0
M17 56 86 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=19140 $dt=0
M18 137 24 89 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=19150 $dt=0
M19 5 25 137 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=19150 $dt=0
M20 57 89 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=19140 $dt=0
M21 5 92 58 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=19140 $dt=0
M22 140 28 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=19150 $dt=0
M23 92 30 140 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=19150 $dt=0
M24 6 62 33 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M25 106 3 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=950 $Y=14910 $dt=1
M26 105 33 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=800 $dt=1
M27 149 51 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M28 41 2 3 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=1880 $Y=14910 $dt=1
M29 4 41 33 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=800 $dt=1
M30 106 64 41 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=2810 $Y=14910 $dt=1
M31 105 63 4 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=800 $dt=1
M32 6 2 64 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=3740 $Y=14910 $dt=1
M33 6 41 63 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=800 $dt=1
M34 108 1 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=14910 $dt=1
M35 66 1 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=20590 $dt=1
M36 6 7 66 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=20590 $dt=1
M37 42 7 1 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=14910 $dt=1
M38 67 42 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=800 $dt=1
M39 108 65 42 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=14910 $dt=1
M40 8 67 107 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=800 $dt=1
M41 6 7 65 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=14910 $dt=1
M42 51 66 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=8230 $Y=20400 $dt=1
M43 34 42 8 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=800 $dt=1
M44 6 34 107 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=800 $dt=1
M45 69 43 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M46 110 9 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M47 70 9 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=20590 $dt=1
M48 6 10 70 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=20590 $dt=1
M49 11 69 111 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M50 43 10 9 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M51 35 43 11 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M52 110 68 43 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M53 6 35 111 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M54 6 10 68 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M55 52 70 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17020 $Y=20400 $dt=1
M56 72 44 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M57 113 12 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M58 73 12 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=20590 $dt=1
M59 14 72 114 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M60 6 13 73 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=20590 $dt=1
M61 44 13 12 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M62 36 44 14 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M63 113 71 44 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M64 6 36 114 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M65 6 13 71 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M66 53 73 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22610 $Y=20400 $dt=1
M67 74 45 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M68 16 74 116 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M69 37 45 16 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M70 6 37 116 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M71 6 78 37 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M72 6 80 54 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27560 $Y=20400 $dt=1
M73 79 15 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M74 159 55 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M75 45 79 127 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M76 17 15 45 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M77 80 15 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29780 $Y=20590 $dt=1
M78 6 17 80 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30190 $Y=20590 $dt=1
M79 6 17 127 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M80 129 18 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M81 82 18 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=20590 $dt=1
M82 6 19 82 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=20590 $dt=1
M83 46 19 18 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M84 83 46 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M85 129 81 46 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M86 20 83 131 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M87 6 19 81 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M88 55 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=34920 $Y=20400 $dt=1
M89 38 46 20 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M90 6 38 131 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M91 85 47 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M92 132 21 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M93 86 21 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=20590 $dt=1
M94 6 22 86 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=20590 $dt=1
M95 23 85 133 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M96 47 22 21 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M97 39 47 23 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M98 132 84 47 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M99 6 39 133 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M100 6 22 84 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M101 56 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=43710 $Y=20400 $dt=1
M102 88 48 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M103 135 24 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M104 89 24 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=20590 $dt=1
M105 27 88 136 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M106 6 25 89 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=20590 $dt=1
M107 48 25 24 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M108 40 48 27 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=48010 $Y=800 $dt=1
M109 135 87 48 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M110 6 40 136 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=48940 $Y=800 $dt=1
M111 6 25 87 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M112 57 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=49300 $Y=20400 $dt=1
M113 138 50 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=50070 $Y=800 $dt=1
M114 26 49 50 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=51000 $Y=800 $dt=1
M115 138 90 26 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=51930 $Y=800 $dt=1
M116 6 49 90 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=52860 $Y=800 $dt=1
M117 6 92 58 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=54210 $Y=20400 $dt=1
M118 91 28 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M119 49 91 139 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M120 164 94 50 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=55830 $Y=11700 $dt=1
M121 6 93 164 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56040 $Y=11700 $dt=1
M122 30 28 49 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M123 92 28 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=20590 $dt=1
M124 6 30 92 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=20590 $dt=1
M125 6 93 163 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56970 $Y=11700 $dt=1
M126 6 30 139 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M127 163 94 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57380 $Y=11700 $dt=1
M128 29 32 163 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57790 $Y=11700 $dt=1
M129 163 31 29 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=58200 $Y=11700 $dt=1
M130 6 31 93 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=59130 $Y=11700 $dt=1
M131 6 32 94 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=60060 $Y=11700 $dt=1
.ends WallaceFinalAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceProject                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceProject 166 165 164 163 162 161 160 159 158 168
+ 169 170 171 172 173 174 93 167 201 200
+ 199 198 197 144 156 154 152 150 206 204
+ 205 203 202 96
** N=656 EP=34 FDC=1660
X0 1 M2_M1_CDNS_765593305580 $T=53500 200590 0 0 $X=53420 $Y=200340
X1 2 M2_M1_CDNS_765593305580 $T=54550 200840 0 0 $X=54470 $Y=200590
X2 3 M2_M1_CDNS_765593305580 $T=73770 191330 0 0 $X=73690 $Y=191080
X3 4 M4_M3_CDNS_765593305581 $T=58900 209500 0 0 $X=58820 $Y=209250
X4 3 M4_M3_CDNS_765593305581 $T=73770 191330 0 0 $X=73690 $Y=191080
X5 1 M3_M2_CDNS_765593305582 $T=53500 200590 0 0 $X=53420 $Y=200340
X6 2 M3_M2_CDNS_765593305582 $T=54550 200840 0 0 $X=54470 $Y=200590
X7 3 M3_M2_CDNS_765593305582 $T=73770 191330 0 0 $X=73690 $Y=191080
X8 5 M2_M1_CDNS_765593305583 $T=35620 163120 0 0 $X=35490 $Y=163040
X9 6 M2_M1_CDNS_765593305583 $T=35930 184200 0 0 $X=35800 $Y=184120
X10 6 M2_M1_CDNS_765593305583 $T=35930 200680 0 0 $X=35800 $Y=200600
X11 7 M2_M1_CDNS_765593305583 $T=36240 154720 0 0 $X=36110 $Y=154640
X12 8 M2_M1_CDNS_765593305583 $T=36550 160830 0 0 $X=36420 $Y=160750
X13 6 M2_M1_CDNS_765593305583 $T=37700 200680 0 0 $X=37570 $Y=200600
X14 9 M2_M1_CDNS_765593305583 $T=38830 161500 0 0 $X=38700 $Y=161420
X15 10 M2_M1_CDNS_765593305583 $T=38870 194470 0 0 $X=38740 $Y=194390
X16 11 M2_M1_CDNS_765593305583 $T=38940 201000 0 0 $X=38810 $Y=200920
X17 7 M2_M1_CDNS_765593305583 $T=39480 154720 0 0 $X=39350 $Y=154640
X18 12 M2_M1_CDNS_765593305583 $T=39480 178900 0 0 $X=39350 $Y=178820
X19 13 M2_M1_CDNS_765593305583 $T=40320 179250 0 0 $X=40190 $Y=179170
X20 14 M2_M1_CDNS_765593305583 $T=40430 161950 0 0 $X=40300 $Y=161870
X21 15 M2_M1_CDNS_765593305583 $T=40520 186280 0 0 $X=40390 $Y=186200
X22 16 M2_M1_CDNS_765593305583 $T=42200 171410 0 0 $X=42070 $Y=171330
X23 17 M2_M1_CDNS_765593305583 $T=42230 193320 0 0 $X=42100 $Y=193240
X24 8 M2_M1_CDNS_765593305583 $T=42850 160830 0 0 $X=42720 $Y=160750
X25 18 M2_M1_CDNS_765593305583 $T=42860 171770 0 0 $X=42730 $Y=171690
X26 19 M2_M1_CDNS_765593305583 $T=43970 180030 0 0 $X=43840 $Y=179950
X27 20 M2_M1_CDNS_765593305583 $T=44740 169870 0 0 $X=44610 $Y=169790
X28 21 M2_M1_CDNS_765593305583 $T=45110 178650 0 0 $X=44980 $Y=178570
X29 22 M2_M1_CDNS_765593305583 $T=45110 190160 0 0 $X=44980 $Y=190080
X30 23 M2_M1_CDNS_765593305583 $T=45550 171360 0 0 $X=45420 $Y=171280
X31 5 M2_M1_CDNS_765593305583 $T=46030 163120 0 0 $X=45900 $Y=163040
X32 24 M2_M1_CDNS_765593305583 $T=46250 169090 0 0 $X=46120 $Y=169010
X33 25 M2_M1_CDNS_765593305583 $T=46270 189090 0 0 $X=46140 $Y=189010
X34 26 M2_M1_CDNS_765593305583 $T=46340 161650 0 0 $X=46210 $Y=161570
X35 27 M2_M1_CDNS_765593305583 $T=47120 186790 0 0 $X=46990 $Y=186710
X36 28 M2_M1_CDNS_765593305583 $T=50150 194020 0 0 $X=50020 $Y=193940
X37 10 M2_M1_CDNS_765593305583 $T=50170 169440 0 0 $X=50040 $Y=169360
X38 29 M2_M1_CDNS_765593305583 $T=50210 163570 0 0 $X=50080 $Y=163490
X39 30 M2_M1_CDNS_765593305583 $T=50210 172170 0 0 $X=50080 $Y=172090
X40 26 M2_M1_CDNS_765593305583 $T=50890 161650 0 0 $X=50760 $Y=161570
X41 31 M2_M1_CDNS_765593305583 $T=50890 188800 0 0 $X=50760 $Y=188720
X42 32 M2_M1_CDNS_765593305583 $T=51310 189500 0 0 $X=51180 $Y=189420
X43 33 M2_M1_CDNS_765593305583 $T=51480 200920 0 0 $X=51350 $Y=200840
X44 3 M2_M1_CDNS_765593305583 $T=51860 186960 0 0 $X=51730 $Y=186880
X45 34 M2_M1_CDNS_765593305583 $T=53210 177850 0 0 $X=53080 $Y=177770
X46 35 M2_M1_CDNS_765593305583 $T=54550 161600 0 0 $X=54420 $Y=161520
X47 36 M2_M1_CDNS_765593305583 $T=54580 170800 0 0 $X=54450 $Y=170720
X48 37 M2_M1_CDNS_765593305583 $T=55280 171060 0 0 $X=55150 $Y=170980
X49 12 M2_M1_CDNS_765593305583 $T=56450 178900 0 0 $X=56320 $Y=178820
X50 38 M2_M1_CDNS_765593305583 $T=56450 192730 0 0 $X=56320 $Y=192650
X51 29 M2_M1_CDNS_765593305583 $T=56870 161900 0 0 $X=56740 $Y=161820
X52 37 M2_M1_CDNS_765593305583 $T=59240 171060 0 0 $X=59110 $Y=170980
X53 37 M2_M1_CDNS_765593305583 $T=59240 171660 0 0 $X=59110 $Y=171580
X54 17 M2_M1_CDNS_765593305583 $T=60710 191070 0 0 $X=60580 $Y=190990
X55 39 M2_M1_CDNS_765593305583 $T=61490 169570 0 0 $X=61360 $Y=169490
X56 40 M2_M1_CDNS_765593305583 $T=61490 186850 0 0 $X=61360 $Y=186770
X57 41 M2_M1_CDNS_765593305583 $T=62210 154420 0 0 $X=62080 $Y=154340
X58 35 M2_M1_CDNS_765593305583 $T=62230 161600 0 0 $X=62100 $Y=161520
X59 42 M2_M1_CDNS_765593305583 $T=62230 187080 0 0 $X=62100 $Y=187000
X60 43 M2_M1_CDNS_765593305583 $T=64550 161600 0 0 $X=64420 $Y=161520
X61 44 M2_M1_CDNS_765593305583 $T=64550 168970 0 0 $X=64420 $Y=168890
X62 45 M2_M1_CDNS_765593305583 $T=64550 178900 0 0 $X=64420 $Y=178820
X63 46 M2_M1_CDNS_765593305583 $T=65890 162940 0 0 $X=65760 $Y=162860
X64 47 M2_M1_CDNS_765593305583 $T=65890 171430 0 0 $X=65760 $Y=171350
X65 48 M2_M1_CDNS_765593305583 $T=65890 179600 0 0 $X=65760 $Y=179520
X66 33 M2_M1_CDNS_765593305583 $T=66830 188900 0 0 $X=66700 $Y=188820
X67 49 M2_M1_CDNS_765593305583 $T=67750 190250 0 0 $X=67620 $Y=190170
X68 43 M2_M1_CDNS_765593305583 $T=68210 161600 0 0 $X=68080 $Y=161520
X69 50 M2_M1_CDNS_765593305583 $T=68210 187730 0 0 $X=68080 $Y=187650
X70 51 M2_M1_CDNS_765593305583 $T=68950 162590 0 0 $X=68820 $Y=162510
X71 52 M2_M1_CDNS_765593305583 $T=68950 186750 0 0 $X=68820 $Y=186670
X72 24 M2_M1_CDNS_765593305583 $T=70970 191030 0 0 $X=70840 $Y=190950
X73 46 M2_M1_CDNS_765593305583 $T=71620 162940 0 0 $X=71490 $Y=162860
X74 25 M2_M1_CDNS_765593305583 $T=71750 186460 0 0 $X=71620 $Y=186380
X75 28 M2_M1_CDNS_765593305583 $T=72150 186680 0 0 $X=72020 $Y=186600
X76 53 M2_M1_CDNS_765593305583 $T=72830 170470 0 0 $X=72700 $Y=170390
X77 47 M2_M1_CDNS_765593305583 $T=73570 171430 0 0 $X=73440 $Y=171350
X78 54 M2_M1_CDNS_765593305583 $T=75890 161600 0 0 $X=75760 $Y=161520
X79 55 M2_M1_CDNS_765593305583 $T=75890 170880 0 0 $X=75760 $Y=170800
X80 56 M2_M1_CDNS_765593305583 $T=77230 161900 0 0 $X=77100 $Y=161820
X81 57 M2_M1_CDNS_765593305583 $T=77530 188080 0 0 $X=77400 $Y=188000
X82 54 M2_M1_CDNS_765593305583 $T=79550 161600 0 0 $X=79420 $Y=161520
X83 58 M2_M1_CDNS_765593305583 $T=79550 178900 0 0 $X=79420 $Y=178820
X84 59 M2_M1_CDNS_765593305583 $T=80240 191050 0 0 $X=80110 $Y=190970
X85 60 M2_M1_CDNS_765593305583 $T=80290 161160 0 0 $X=80160 $Y=161080
X86 30 M2_M1_CDNS_765593305583 $T=80290 169870 0 0 $X=80160 $Y=169790
X87 61 M2_M1_CDNS_765593305583 $T=80290 188490 0 0 $X=80160 $Y=188410
X88 62 M2_M1_CDNS_765593305583 $T=80570 189620 0 0 $X=80440 $Y=189540
X89 63 M2_M1_CDNS_765593305583 $T=82800 189650 0 0 $X=82670 $Y=189570
X90 64 M2_M1_CDNS_765593305583 $T=84170 170170 0 0 $X=84040 $Y=170090
X91 65 M2_M1_CDNS_765593305583 $T=84170 178140 0 0 $X=84040 $Y=178060
X92 66 M2_M1_CDNS_765593305583 $T=84300 154200 0 0 $X=84170 $Y=154120
X93 67 M2_M1_CDNS_765593305583 $T=84910 179770 0 0 $X=84780 $Y=179690
X94 68 M2_M1_CDNS_765593305583 $T=84920 188870 0 0 $X=84790 $Y=188790
X95 40 M2_M1_CDNS_765593305583 $T=85640 189410 0 0 $X=85510 $Y=189330
X96 69 M2_M1_CDNS_765593305583 $T=87590 186550 0 0 $X=87460 $Y=186470
X97 61 M2_M1_CDNS_765593305583 $T=88020 188490 0 0 $X=87890 $Y=188410
X98 70 M2_M1_CDNS_765593305583 $T=88260 171660 0 0 $X=88130 $Y=171580
X99 71 M2_M1_CDNS_765593305583 $T=90090 186600 0 0 $X=89960 $Y=186520
X100 72 M2_M1_CDNS_765593305583 $T=90500 188430 0 0 $X=90370 $Y=188350
X101 72 M2_M1_CDNS_765593305583 $T=90500 189690 0 0 $X=90370 $Y=189610
X102 73 M2_M1_CDNS_765593305583 $T=91320 186600 0 0 $X=91190 $Y=186520
X103 74 M2_M1_CDNS_765593305583 $T=91570 163270 0 0 $X=91440 $Y=163190
X104 75 M2_M1_CDNS_765593305583 $T=91610 161180 0 0 $X=91480 $Y=161100
X105 50 M2_M1_CDNS_765593305583 $T=94040 190140 0 0 $X=93910 $Y=190060
X106 76 M2_M1_CDNS_765593305583 $T=94390 190970 0 0 $X=94260 $Y=190890
X107 77 M2_M1_CDNS_765593305583 $T=95520 170420 0 0 $X=95390 $Y=170340
X108 73 M2_M1_CDNS_765593305583 $T=98230 186600 0 0 $X=98100 $Y=186520
X109 5 M3_M2_CDNS_765593305584 $T=35620 163120 0 0 $X=35490 $Y=162750
X110 6 M3_M2_CDNS_765593305584 $T=35930 184200 0 0 $X=35800 $Y=183830
X111 12 M3_M2_CDNS_765593305584 $T=39480 178900 0 0 $X=39350 $Y=178530
X112 78 M3_M2_CDNS_765593305584 $T=39970 179890 0 0 $X=39840 $Y=179520
X113 13 M3_M2_CDNS_765593305584 $T=40320 179250 0 0 $X=40190 $Y=178880
X114 16 M3_M2_CDNS_765593305584 $T=42200 171410 0 0 $X=42070 $Y=171040
X115 36 M3_M2_CDNS_765593305584 $T=42900 200500 0 0 $X=42770 $Y=200130
X116 79 M3_M2_CDNS_765593305584 $T=45110 201840 0 0 $X=44980 $Y=201470
X117 24 M3_M2_CDNS_765593305584 $T=46250 169090 0 0 $X=46120 $Y=168720
X118 80 M3_M2_CDNS_765593305584 $T=46270 179600 0 0 $X=46140 $Y=179230
X119 81 M3_M2_CDNS_765593305584 $T=46270 201250 0 0 $X=46140 $Y=200880
X120 27 M3_M2_CDNS_765593305584 $T=47120 186790 0 0 $X=46990 $Y=186420
X121 82 M3_M2_CDNS_765593305584 $T=50150 201310 0 0 $X=50020 $Y=200940
X122 33 M3_M2_CDNS_765593305584 $T=51480 200920 0 0 $X=51350 $Y=200550
X123 39 M3_M2_CDNS_765593305584 $T=54200 207730 0 0 $X=54070 $Y=207360
X124 3 M3_M2_CDNS_765593305584 $T=55250 191340 0 0 $X=55120 $Y=190970
X125 83 M3_M2_CDNS_765593305584 $T=55950 186300 0 0 $X=55820 $Y=185930
X126 84 M3_M2_CDNS_765593305584 $T=56870 188050 0 0 $X=56740 $Y=187680
X127 85 M3_M2_CDNS_765593305584 $T=57590 186350 0 0 $X=57460 $Y=185980
X128 1 M3_M2_CDNS_765593305584 $T=57610 178190 0 0 $X=57480 $Y=177820
X129 86 M3_M2_CDNS_765593305584 $T=61520 191010 0 0 $X=61390 $Y=190640
X130 87 M3_M2_CDNS_765593305584 $T=61840 177950 0 0 $X=61710 $Y=177580
X131 82 M3_M2_CDNS_765593305584 $T=62320 191010 0 0 $X=62190 $Y=190640
X132 50 M3_M2_CDNS_765593305584 $T=68210 187730 0 0 $X=68080 $Y=187360
X133 20 M3_M2_CDNS_765593305584 $T=68950 169520 0 0 $X=68820 $Y=169150
X134 24 M3_M2_CDNS_765593305584 $T=70970 191030 0 0 $X=70840 $Y=190660
X135 88 M3_M2_CDNS_765593305584 $T=72950 189120 0 0 $X=72820 $Y=188750
X136 48 M3_M2_CDNS_765593305584 $T=73180 177950 0 0 $X=73050 $Y=177580
X137 89 M3_M2_CDNS_765593305584 $T=73260 186550 0 0 $X=73130 $Y=186180
X138 90 M3_M2_CDNS_765593305584 $T=75390 187080 0 0 $X=75260 $Y=186710
X139 91 M3_M2_CDNS_765593305584 $T=79550 189730 0 0 $X=79420 $Y=189360
X140 64 M3_M2_CDNS_765593305584 $T=84170 170170 0 0 $X=84040 $Y=169800
X141 92 M3_M2_CDNS_765593305584 $T=91630 178250 0 0 $X=91500 $Y=177880
X142 50 M3_M2_CDNS_765593305584 $T=94040 190140 0 0 $X=93910 $Y=189770
X143 93 M3_M2_CDNS_765593305585 $T=36870 154210 0 0 $X=36790 $Y=153960
X144 94 M3_M2_CDNS_765593305585 $T=39090 200490 0 0 $X=39010 $Y=200240
X145 95 M3_M2_CDNS_765593305585 $T=43880 210410 0 0 $X=43800 $Y=210160
X146 93 M3_M2_CDNS_765593305585 $T=48210 153790 0 0 $X=48130 $Y=153540
X147 96 M3_M2_CDNS_765593305585 $T=53980 160640 0 0 $X=53900 $Y=160390
X148 41 M3_M2_CDNS_765593305585 $T=59140 149330 0 0 $X=59060 $Y=149080
X149 93 M3_M2_CDNS_765593305585 $T=59550 153740 0 0 $X=59470 $Y=153490
X150 2 M3_M2_CDNS_765593305585 $T=61490 178760 0 0 $X=61410 $Y=178510
X151 96 M3_M2_CDNS_765593305585 $T=65090 160640 0 0 $X=65010 $Y=160390
X152 93 M3_M2_CDNS_765593305585 $T=70770 153700 0 0 $X=70690 $Y=153450
X153 97 M3_M2_CDNS_765593305585 $T=71450 149330 0 0 $X=71370 $Y=149080
X154 96 M3_M2_CDNS_765593305585 $T=76650 169330 0 0 $X=76570 $Y=169080
X155 93 M3_M2_CDNS_765593305585 $T=82230 153680 0 0 $X=82150 $Y=153430
X156 96 M3_M2_CDNS_765593305585 $T=87810 169220 0 0 $X=87730 $Y=168970
X157 93 M3_M2_CDNS_765593305585 $T=93570 153650 0 0 $X=93490 $Y=153400
X158 93 M3_M2_CDNS_765593305585 $T=95590 138740 0 180 $X=95510 $Y=138490
X159 5 M2_M1_CDNS_765593305586 $T=35620 207840 0 0 $X=35540 $Y=207710
X160 7 M2_M1_CDNS_765593305586 $T=36240 193000 0 0 $X=36160 $Y=192870
X161 5 M2_M1_CDNS_765593305586 $T=37600 210470 0 0 $X=37520 $Y=210340
X162 88 M2_M1_CDNS_765593305586 $T=37880 178170 0 0 $X=37800 $Y=178040
X163 86 M2_M1_CDNS_765593305586 $T=38450 201870 0 0 $X=38370 $Y=201740
X164 98 M2_M1_CDNS_765593305586 $T=38810 170080 0 0 $X=38730 $Y=169950
X165 99 M2_M1_CDNS_765593305586 $T=38830 187050 0 0 $X=38750 $Y=186920
X166 100 M2_M1_CDNS_765593305586 $T=38870 187540 0 0 $X=38790 $Y=187410
X167 87 M2_M1_CDNS_765593305586 $T=39150 180820 0 0 $X=39070 $Y=180690
X168 7 M2_M1_CDNS_765593305586 $T=39190 193000 0 0 $X=39110 $Y=192870
X169 101 M2_M1_CDNS_765593305586 $T=39480 194520 0 0 $X=39400 $Y=194390
X170 51 M2_M1_CDNS_765593305586 $T=39530 162590 0 0 $X=39450 $Y=162460
X171 96 M2_M1_CDNS_765593305586 $T=39560 210360 0 0 $X=39480 $Y=210230
X172 101 M2_M1_CDNS_765593305586 $T=39860 200520 0 0 $X=39780 $Y=200390
X173 78 M2_M1_CDNS_765593305586 $T=39970 179890 0 0 $X=39890 $Y=179760
X174 49 M2_M1_CDNS_765593305586 $T=40830 171740 0 0 $X=40750 $Y=171610
X175 20 M2_M1_CDNS_765593305586 $T=41870 163060 0 0 $X=41790 $Y=162930
X176 96 M2_M1_CDNS_765593305586 $T=42470 210800 0 0 $X=42390 $Y=210670
X177 18 M2_M1_CDNS_765593305586 $T=42860 186180 0 0 $X=42780 $Y=186050
X178 18 M2_M1_CDNS_765593305586 $T=42860 194640 0 0 $X=42780 $Y=194510
X179 36 M2_M1_CDNS_765593305586 $T=42900 200500 0 0 $X=42820 $Y=200370
X180 53 M2_M1_CDNS_765593305586 $T=43210 170470 0 0 $X=43130 $Y=170340
X181 62 M2_M1_CDNS_765593305586 $T=44650 186080 0 0 $X=44570 $Y=185950
X182 102 M2_M1_CDNS_765593305586 $T=44700 186580 0 0 $X=44620 $Y=186450
X183 20 M2_M1_CDNS_765593305586 $T=44740 168980 0 0 $X=44660 $Y=168850
X184 79 M2_M1_CDNS_765593305586 $T=45110 201840 0 0 $X=45030 $Y=201710
X185 93 M2_M1_CDNS_765593305586 $T=45220 210430 0 0 $X=45140 $Y=210300
X186 59 M2_M1_CDNS_765593305586 $T=45530 187610 0 0 $X=45450 $Y=187480
X187 80 M2_M1_CDNS_765593305586 $T=46270 179600 0 0 $X=46190 $Y=179470
X188 81 M2_M1_CDNS_765593305586 $T=46270 201250 0 0 $X=46190 $Y=201120
X189 103 M2_M1_CDNS_765593305586 $T=46870 210480 0 0 $X=46790 $Y=210350
X190 28 M2_M1_CDNS_765593305586 $T=47730 186910 0 0 $X=47650 $Y=186780
X191 28 M2_M1_CDNS_765593305586 $T=47730 194020 0 0 $X=47650 $Y=193890
X192 93 M2_M1_CDNS_765593305586 $T=48140 210720 0 0 $X=48060 $Y=210590
X193 104 M2_M1_CDNS_765593305586 $T=48860 186230 0 0 $X=48780 $Y=186100
X194 95 M2_M1_CDNS_765593305586 $T=49200 172030 0 0 $X=49120 $Y=171900
X195 105 M2_M1_CDNS_765593305586 $T=49540 210490 0 0 $X=49460 $Y=210360
X196 103 M2_M1_CDNS_765593305586 $T=50150 160980 0 0 $X=50070 $Y=160850
X197 82 M2_M1_CDNS_765593305586 $T=50150 201310 0 0 $X=50070 $Y=201180
X198 96 M2_M1_CDNS_765593305586 $T=50900 210460 0 0 $X=50820 $Y=210330
X199 96 M2_M1_CDNS_765593305586 $T=51730 210520 0 0 $X=51650 $Y=210390
X200 106 M2_M1_CDNS_765593305586 $T=52160 180360 0 0 $X=52080 $Y=180230
X201 107 M2_M1_CDNS_765593305586 $T=52210 186080 0 0 $X=52130 $Y=185950
X202 108 M2_M1_CDNS_765593305586 $T=52520 210480 0 0 $X=52440 $Y=210350
X203 60 M2_M1_CDNS_765593305586 $T=52690 169020 0 0 $X=52610 $Y=168890
X204 60 M2_M1_CDNS_765593305586 $T=54180 161160 0 0 $X=54100 $Y=161030
X205 60 M2_M1_CDNS_765593305586 $T=54180 165330 0 0 $X=54100 $Y=165200
X206 39 M2_M1_CDNS_765593305586 $T=55230 210480 0 0 $X=55150 $Y=210350
X207 83 M2_M1_CDNS_765593305586 $T=55950 186230 0 0 $X=55870 $Y=186100
X208 109 M2_M1_CDNS_765593305586 $T=56450 200950 0 0 $X=56370 $Y=200820
X209 93 M2_M1_CDNS_765593305586 $T=56570 210480 0 0 $X=56490 $Y=210350
X210 63 M2_M1_CDNS_765593305586 $T=56860 180370 0 0 $X=56780 $Y=180240
X211 84 M2_M1_CDNS_765593305586 $T=56870 188050 0 0 $X=56790 $Y=187920
X212 64 M2_M1_CDNS_765593305586 $T=56940 181050 0 0 $X=56860 $Y=180920
X213 85 M2_M1_CDNS_765593305586 $T=57590 186230 0 0 $X=57510 $Y=186100
X214 1 M2_M1_CDNS_765593305586 $T=57610 178190 0 0 $X=57530 $Y=178060
X215 105 M2_M1_CDNS_765593305586 $T=57700 162210 0 0 $X=57620 $Y=162080
X216 4 M2_M1_CDNS_765593305586 $T=58210 210480 0 0 $X=58130 $Y=210350
X217 65 M2_M1_CDNS_765593305586 $T=58360 177710 0 0 $X=58280 $Y=177580
X218 110 M2_M1_CDNS_765593305586 $T=58700 201250 0 0 $X=58620 $Y=201120
X219 111 M2_M1_CDNS_765593305586 $T=59000 193970 0 0 $X=58920 $Y=193840
X220 93 M2_M1_CDNS_765593305586 $T=59490 210790 0 0 $X=59410 $Y=210660
X221 14 M2_M1_CDNS_765593305586 $T=60200 186560 0 0 $X=60120 $Y=186430
X222 81 M2_M1_CDNS_765593305586 $T=60650 186550 0 0 $X=60570 $Y=186420
X223 4 M2_M1_CDNS_765593305586 $T=61490 162160 0 0 $X=61410 $Y=162030
X224 86 M2_M1_CDNS_765593305586 $T=61520 191010 0 0 $X=61440 $Y=190880
X225 87 M2_M1_CDNS_765593305586 $T=61840 177950 0 0 $X=61760 $Y=177820
X226 37 M2_M1_CDNS_765593305586 $T=62230 171360 0 0 $X=62150 $Y=171230
X227 82 M2_M1_CDNS_765593305586 $T=62320 191010 0 0 $X=62240 $Y=190880
X228 112 M2_M1_CDNS_765593305586 $T=62650 188450 0 0 $X=62570 $Y=188320
X229 110 M2_M1_CDNS_765593305586 $T=62720 191010 0 0 $X=62640 $Y=190880
X230 98 M2_M1_CDNS_765593305586 $T=62980 190210 0 0 $X=62900 $Y=190080
X231 80 M2_M1_CDNS_765593305586 $T=63540 186400 0 0 $X=63460 $Y=186270
X232 106 M2_M1_CDNS_765593305586 $T=63920 187450 0 0 $X=63840 $Y=187320
X233 9 M2_M1_CDNS_765593305586 $T=65000 188900 0 0 $X=64920 $Y=188770
X234 11 M2_M1_CDNS_765593305586 $T=66120 189270 0 0 $X=66040 $Y=189140
X235 44 M2_M1_CDNS_765593305586 $T=66900 168970 0 0 $X=66820 $Y=168840
X236 109 M2_M1_CDNS_765593305586 $T=67350 188950 0 0 $X=67270 $Y=188820
X237 57 M2_M1_CDNS_765593305586 $T=67790 188080 0 0 $X=67710 $Y=187950
X238 21 M2_M1_CDNS_765593305586 $T=68140 190600 0 0 $X=68060 $Y=190470
X239 45 M2_M1_CDNS_765593305586 $T=68210 178900 0 0 $X=68130 $Y=178770
X240 16 M2_M1_CDNS_765593305586 $T=68610 178140 0 0 $X=68530 $Y=178010
X241 20 M2_M1_CDNS_765593305586 $T=68950 169520 0 0 $X=68870 $Y=169390
X242 94 M2_M1_CDNS_765593305586 $T=70040 186090 0 0 $X=69960 $Y=185960
X243 23 M2_M1_CDNS_765593305586 $T=71980 162150 0 0 $X=71900 $Y=162020
X244 111 M2_M1_CDNS_765593305586 $T=72550 190420 0 0 $X=72470 $Y=190290
X245 19 M2_M1_CDNS_765593305586 $T=72830 179740 0 0 $X=72750 $Y=179610
X246 88 M2_M1_CDNS_765593305586 $T=72950 189120 0 0 $X=72870 $Y=188990
X247 48 M2_M1_CDNS_765593305586 $T=73180 177950 0 0 $X=73100 $Y=177820
X248 89 M2_M1_CDNS_765593305586 $T=73260 186550 0 0 $X=73180 $Y=186420
X249 27 M2_M1_CDNS_765593305586 $T=73340 189950 0 0 $X=73260 $Y=189820
X250 113 M2_M1_CDNS_765593305586 $T=75110 189850 0 0 $X=75030 $Y=189720
X251 90 M2_M1_CDNS_765593305586 $T=75390 187080 0 0 $X=75310 $Y=186950
X252 6 M2_M1_CDNS_765593305586 $T=75810 186640 0 0 $X=75730 $Y=186510
X253 58 M2_M1_CDNS_765593305586 $T=75890 178900 0 0 $X=75810 $Y=178770
X254 22 M2_M1_CDNS_765593305586 $T=76210 186310 0 0 $X=76130 $Y=186180
X255 32 M2_M1_CDNS_765593305586 $T=76610 189710 0 0 $X=76530 $Y=189580
X256 38 M2_M1_CDNS_765593305586 $T=77010 186270 0 0 $X=76930 $Y=186140
X257 114 M2_M1_CDNS_765593305586 $T=77230 171250 0 0 $X=77150 $Y=171120
X258 67 M2_M1_CDNS_765593305586 $T=77230 179770 0 0 $X=77150 $Y=179640
X259 78 M2_M1_CDNS_765593305586 $T=77410 188450 0 0 $X=77330 $Y=188320
X260 102 M2_M1_CDNS_765593305586 $T=77810 189900 0 0 $X=77730 $Y=189770
X261 107 M2_M1_CDNS_765593305586 $T=78220 190490 0 0 $X=78140 $Y=190360
X262 83 M2_M1_CDNS_765593305586 $T=78600 191010 0 0 $X=78520 $Y=190880
X263 84 M2_M1_CDNS_765593305586 $T=78690 189850 0 0 $X=78610 $Y=189720
X264 55 M2_M1_CDNS_765593305586 $T=79550 170880 0 0 $X=79470 $Y=170750
X265 91 M2_M1_CDNS_765593305586 $T=79550 189730 0 0 $X=79470 $Y=189600
X266 115 M2_M1_CDNS_765593305586 $T=79570 153500 0 0 $X=79490 $Y=153370
X267 104 M2_M1_CDNS_765593305586 $T=79890 190750 0 0 $X=79810 $Y=190620
X268 34 M2_M1_CDNS_765593305586 $T=80290 178350 0 0 $X=80210 $Y=178220
X269 61 M2_M1_CDNS_765593305586 $T=80290 186790 0 0 $X=80210 $Y=186660
X270 13 M2_M1_CDNS_765593305586 $T=82110 190200 0 0 $X=82030 $Y=190070
X271 31 M2_M1_CDNS_765593305586 $T=82890 191000 0 0 $X=82810 $Y=190870
X272 85 M2_M1_CDNS_765593305586 $T=83150 190000 0 0 $X=83070 $Y=189870
X273 92 M2_M1_CDNS_765593305586 $T=83710 190340 0 0 $X=83630 $Y=190210
X274 116 M2_M1_CDNS_765593305586 $T=84170 186790 0 0 $X=84090 $Y=186660
X275 56 M2_M1_CDNS_765593305586 $T=84190 161900 0 0 $X=84110 $Y=161770
X276 117 M2_M1_CDNS_765593305586 $T=84840 153500 0 0 $X=84760 $Y=153370
X277 114 M2_M1_CDNS_765593305586 $T=84910 171250 0 0 $X=84830 $Y=171120
X278 68 M2_M1_CDNS_765593305586 $T=84920 187190 0 0 $X=84840 $Y=187060
X279 75 M2_M1_CDNS_765593305586 $T=87230 161180 0 0 $X=87150 $Y=161050
X280 70 M2_M1_CDNS_765593305586 $T=87230 171660 0 0 $X=87150 $Y=171530
X281 118 M2_M1_CDNS_765593305586 $T=87230 178550 0 0 $X=87150 $Y=178420
X282 52 M2_M1_CDNS_765593305586 $T=87230 189630 0 0 $X=87150 $Y=189500
X283 113 M2_M1_CDNS_765593305586 $T=87620 191030 0 0 $X=87540 $Y=190900
X284 61 M2_M1_CDNS_765593305586 $T=88020 189460 0 0 $X=87940 $Y=189330
X285 116 M2_M1_CDNS_765593305586 $T=88410 190610 0 0 $X=88330 $Y=190480
X286 119 M2_M1_CDNS_765593305586 $T=90480 169080 0 0 $X=90400 $Y=168950
X287 119 M2_M1_CDNS_765593305586 $T=90480 171540 0 0 $X=90400 $Y=171410
X288 99 M2_M1_CDNS_765593305586 $T=90620 191090 0 0 $X=90540 $Y=190960
X289 120 M2_M1_CDNS_765593305586 $T=90820 187480 0 0 $X=90740 $Y=187350
X290 118 M2_M1_CDNS_765593305586 $T=90890 178550 0 0 $X=90810 $Y=178420
X291 112 M2_M1_CDNS_765593305586 $T=91420 189850 0 0 $X=91340 $Y=189720
X292 92 M2_M1_CDNS_765593305586 $T=91630 178250 0 0 $X=91550 $Y=178120
X293 90 M2_M1_CDNS_765593305586 $T=92230 189370 0 0 $X=92150 $Y=189240
X294 120 M2_M1_CDNS_765593305586 $T=92620 189600 0 0 $X=92540 $Y=189470
X295 77 M2_M1_CDNS_765593305586 $T=92740 170420 0 0 $X=92660 $Y=170290
X296 69 M2_M1_CDNS_765593305586 $T=93020 190510 0 0 $X=92940 $Y=190380
X297 71 M2_M1_CDNS_765593305586 $T=93410 189290 0 0 $X=93330 $Y=189160
X298 74 M2_M1_CDNS_765593305586 $T=95520 160860 0 0 $X=95440 $Y=160730
X299 76 M2_M1_CDNS_765593305586 $T=95520 188060 0 0 $X=95440 $Y=187930
X300 121 M2_M1_CDNS_765593305586 $T=95530 177680 0 0 $X=95450 $Y=177550
X301 42 M2_M1_CDNS_765593305586 $T=96230 190670 0 0 $X=96150 $Y=190540
X302 89 M2_M1_CDNS_765593305586 $T=97030 190540 0 0 $X=96950 $Y=190410
X303 91 M2_M1_CDNS_765593305586 $T=97430 190230 0 0 $X=97350 $Y=190100
X304 11 M3_M2_CDNS_765593305587 $T=38220 201000 0 0 $X=38090 $Y=200920
X305 98 M3_M2_CDNS_765593305587 $T=38810 172200 0 0 $X=38680 $Y=172120
X306 36 M3_M2_CDNS_765593305587 $T=42900 185000 0 0 $X=42770 $Y=184920
X307 36 M3_M2_CDNS_765593305587 $T=43110 179550 0 0 $X=42980 $Y=179470
X308 103 M3_M2_CDNS_765593305587 $T=43600 185000 0 0 $X=43470 $Y=184920
X309 103 M3_M2_CDNS_765593305587 $T=43600 196610 0 0 $X=43470 $Y=196530
X310 9 M3_M2_CDNS_765593305587 $T=44630 161500 0 0 $X=44500 $Y=161420
X311 19 M3_M2_CDNS_765593305587 $T=45280 180030 0 0 $X=45150 $Y=179950
X312 103 M3_M2_CDNS_765593305587 $T=47510 160980 0 0 $X=47380 $Y=160900
X313 95 M3_M2_CDNS_765593305587 $T=49200 180640 0 0 $X=49070 $Y=180560
X314 12 M3_M2_CDNS_765593305587 $T=49630 178900 0 0 $X=49500 $Y=178820
X315 23 M3_M2_CDNS_765593305587 $T=52770 171360 0 0 $X=52640 $Y=171280
X316 79 M3_M2_CDNS_765593305587 $T=53420 184700 0 0 $X=53290 $Y=184620
X317 15 M3_M2_CDNS_765593305587 $T=53630 188450 0 0 $X=53500 $Y=188370
X318 53 M3_M2_CDNS_765593305587 $T=54580 170470 0 0 $X=54450 $Y=170390
X319 31 M3_M2_CDNS_765593305587 $T=55250 188800 0 0 $X=55120 $Y=188720
X320 53 M3_M2_CDNS_765593305587 $T=56260 170470 0 0 $X=56130 $Y=170390
X321 23 M3_M2_CDNS_765593305587 $T=56630 171360 0 0 $X=56500 $Y=171280
X322 63 M3_M2_CDNS_765593305587 $T=56860 180700 0 0 $X=56730 $Y=180620
X323 20 M3_M2_CDNS_765593305587 $T=57000 170170 0 0 $X=56870 $Y=170090
X324 108 M3_M2_CDNS_765593305587 $T=57350 169570 0 0 $X=57220 $Y=169490
X325 109 M3_M2_CDNS_765593305587 $T=58750 185300 0 0 $X=58620 $Y=185220
X326 14 M3_M2_CDNS_765593305587 $T=60200 180400 0 0 $X=60070 $Y=180320
X327 81 M3_M2_CDNS_765593305587 $T=60650 183850 0 0 $X=60520 $Y=183770
X328 40 M3_M2_CDNS_765593305587 $T=61490 186700 0 0 $X=61360 $Y=186620
X329 80 M3_M2_CDNS_765593305587 $T=63330 186400 0 0 $X=63200 $Y=186320
X330 9 M3_M2_CDNS_765593305587 $T=65000 181400 0 0 $X=64870 $Y=181320
X331 79 M3_M2_CDNS_765593305587 $T=65670 184700 0 0 $X=65540 $Y=184620
X332 79 M3_M2_CDNS_765593305587 $T=65670 191010 0 0 $X=65540 $Y=190930
X333 11 M3_M2_CDNS_765593305587 $T=66120 182800 0 0 $X=65990 $Y=182720
X334 109 M3_M2_CDNS_765593305587 $T=67350 185300 0 0 $X=67220 $Y=185220
X335 49 M3_M2_CDNS_765593305587 $T=67490 190250 0 0 $X=67360 $Y=190170
X336 21 M3_M2_CDNS_765593305587 $T=67930 190600 0 0 $X=67800 $Y=190520
X337 20 M3_M2_CDNS_765593305587 $T=68950 170170 0 0 $X=68820 $Y=170090
X338 94 M3_M2_CDNS_765593305587 $T=70040 183500 0 0 $X=69910 $Y=183420
X339 25 M3_M2_CDNS_765593305587 $T=71750 185000 0 0 $X=71620 $Y=184920
X340 23 M3_M2_CDNS_765593305587 $T=71980 171010 0 0 $X=71850 $Y=170930
X341 28 M3_M2_CDNS_765593305587 $T=72150 185950 0 0 $X=72020 $Y=185870
X342 19 M3_M2_CDNS_765593305587 $T=72830 180030 0 0 $X=72700 $Y=179950
X343 34 M3_M2_CDNS_765593305587 $T=73630 178350 0 0 $X=73500 $Y=178270
X344 6 M3_M2_CDNS_765593305587 $T=75810 184200 0 0 $X=75680 $Y=184120
X345 32 M3_M2_CDNS_765593305587 $T=76610 189500 0 0 $X=76480 $Y=189420
X346 102 M3_M2_CDNS_765593305587 $T=77510 189900 0 0 $X=77380 $Y=189820
X347 83 M3_M2_CDNS_765593305587 $T=77770 185600 0 0 $X=77640 $Y=185520
X348 107 M3_M2_CDNS_765593305587 $T=78220 189850 0 0 $X=78090 $Y=189770
X349 13 M3_M2_CDNS_765593305587 $T=78720 190200 0 0 $X=78590 $Y=190120
X350 91 M3_M2_CDNS_765593305587 $T=82800 187430 0 0 $X=82670 $Y=187350
X351 85 M3_M2_CDNS_765593305587 $T=83150 186700 0 0 $X=83020 $Y=186620
X352 90 M3_M2_CDNS_765593305587 $T=89270 187080 0 0 $X=89140 $Y=187000
X353 122 M2_M1_CDNS_765593305588 $T=36060 153500 0 0 $X=35930 $Y=153370
X354 122 M2_M1_CDNS_765593305588 $T=43210 153500 0 0 $X=43080 $Y=153370
X355 123 M2_M1_CDNS_765593305588 $T=49210 149200 0 0 $X=49080 $Y=149070
X356 123 M2_M1_CDNS_765593305588 $T=49210 153930 0 0 $X=49080 $Y=153800
X357 124 M2_M1_CDNS_765593305588 $T=54550 153500 0 0 $X=54420 $Y=153370
X358 125 M2_M1_CDNS_765593305588 $T=56890 153870 0 0 $X=56760 $Y=153740
X359 108 M2_M1_CDNS_765593305588 $T=57610 169570 0 0 $X=57480 $Y=169440
X360 126 M2_M1_CDNS_765593305588 $T=63660 149840 0 0 $X=63530 $Y=149710
X361 127 M2_M1_CDNS_765593305588 $T=64550 153500 0 0 $X=64420 $Y=153370
X362 79 M2_M1_CDNS_765593305588 $T=66540 191010 0 0 $X=66410 $Y=190880
X363 127 M2_M1_CDNS_765593305588 $T=67160 148490 0 0 $X=67030 $Y=148360
X364 128 M2_M1_CDNS_765593305588 $T=67780 149140 0 0 $X=67650 $Y=149010
X365 97 M2_M1_CDNS_765593305588 $T=73550 154200 0 0 $X=73420 $Y=154070
X366 129 M2_M1_CDNS_765593305588 $T=77230 154200 0 0 $X=77100 $Y=154070
X367 15 M2_M1_CDNS_765593305588 $T=86440 190310 0 0 $X=86310 $Y=190180
X368 130 M2_M1_CDNS_765593305588 $T=90300 149720 0 0 $X=90170 $Y=149590
X369 130 M2_M1_CDNS_765593305588 $T=90960 153490 0 0 $X=90830 $Y=153360
X370 131 M2_M1_CDNS_765593305588 $T=91570 155020 0 0 $X=91440 $Y=154890
X371 10 M3_M2_CDNS_765593305589 $T=37650 169730 0 0 $X=37570 $Y=169600
X372 10 M3_M2_CDNS_765593305589 $T=37650 193960 0 0 $X=37570 $Y=193830
X373 86 M3_M2_CDNS_765593305589 $T=38570 200640 0 0 $X=38490 $Y=200510
X374 86 M3_M2_CDNS_765593305589 $T=38570 201610 0 0 $X=38490 $Y=201480
X375 88 M3_M2_CDNS_765593305589 $T=39000 178170 0 0 $X=38920 $Y=178040
X376 99 M3_M2_CDNS_765593305589 $T=39350 187050 0 0 $X=39270 $Y=186920
X377 49 M3_M2_CDNS_765593305589 $T=40830 172550 0 0 $X=40750 $Y=172420
X378 87 M3_M2_CDNS_765593305589 $T=41330 177500 0 0 $X=41250 $Y=177370
X379 21 M3_M2_CDNS_765593305589 $T=42600 184650 0 0 $X=42520 $Y=184520
X380 62 M3_M2_CDNS_765593305589 $T=44650 185230 0 0 $X=44570 $Y=185100
X381 22 M3_M2_CDNS_765593305589 $T=45350 190160 0 0 $X=45270 $Y=190030
X382 59 M3_M2_CDNS_765593305589 $T=46050 187610 0 0 $X=45970 $Y=187480
X383 103 M3_M2_CDNS_765593305589 $T=47510 178550 0 0 $X=47430 $Y=178420
X384 28 M3_M2_CDNS_765593305589 $T=47730 185950 0 0 $X=47650 $Y=185820
X385 25 M3_M2_CDNS_765593305589 $T=48030 185000 0 0 $X=47950 $Y=184870
X386 25 M3_M2_CDNS_765593305589 $T=48030 186910 0 0 $X=47950 $Y=186780
X387 25 M3_M2_CDNS_765593305589 $T=48030 189090 0 0 $X=47950 $Y=188960
X388 104 M3_M2_CDNS_765593305589 $T=48860 183960 0 0 $X=48780 $Y=183830
X389 107 M3_M2_CDNS_765593305589 $T=52210 183840 0 0 $X=52130 $Y=183710
X390 105 M3_M2_CDNS_765593305589 $T=53150 207870 0 0 $X=53070 $Y=207740
X391 29 M3_M2_CDNS_765593305589 $T=53240 163570 0 0 $X=53160 $Y=163440
X392 79 M3_M2_CDNS_765593305589 $T=53420 186300 0 0 $X=53340 $Y=186170
X393 108 M3_M2_CDNS_765593305589 $T=53890 207420 0 0 $X=53810 $Y=207290
X394 32 M3_M2_CDNS_765593305589 $T=53900 189500 0 0 $X=53820 $Y=189370
X395 3 M3_M2_CDNS_765593305589 $T=54460 187880 0 0 $X=54380 $Y=187750
X396 3 M3_M2_CDNS_765593305589 $T=54460 189220 0 0 $X=54380 $Y=189090
X397 64 M3_M2_CDNS_765593305589 $T=58010 176100 0 0 $X=57930 $Y=175970
X398 65 M3_M2_CDNS_765593305589 $T=58360 175400 0 0 $X=58280 $Y=175270
X399 109 M3_M2_CDNS_765593305589 $T=58750 186300 0 0 $X=58670 $Y=186170
X400 98 M3_M2_CDNS_765593305589 $T=59010 188800 0 0 $X=58930 $Y=188670
X401 27 M3_M2_CDNS_765593305589 $T=63360 189950 0 0 $X=63280 $Y=189820
X402 112 M3_M2_CDNS_765593305589 $T=63730 188450 0 0 $X=63650 $Y=188320
X403 79 M3_M2_CDNS_765593305589 $T=65670 188550 0 0 $X=65590 $Y=188420
X404 33 M3_M2_CDNS_765593305589 $T=66830 183140 0 0 $X=66750 $Y=183010
X405 48 M3_M2_CDNS_765593305589 $T=67770 179600 0 0 $X=67690 $Y=179470
X406 16 M3_M2_CDNS_765593305589 $T=68610 176870 0 0 $X=68530 $Y=176740
X407 23 M3_M2_CDNS_765593305589 $T=71980 162410 0 0 $X=71900 $Y=162280
X408 111 M3_M2_CDNS_765593305589 $T=72550 190680 0 0 $X=72470 $Y=190550
X409 111 M3_M2_CDNS_765593305589 $T=72550 193970 0 0 $X=72470 $Y=193840
X410 113 M3_M2_CDNS_765593305589 $T=75110 190970 0 0 $X=75030 $Y=190840
X411 22 M3_M2_CDNS_765593305589 $T=76210 185600 0 0 $X=76130 $Y=185470
X412 38 M3_M2_CDNS_765593305589 $T=77010 185650 0 0 $X=76930 $Y=185520
X413 78 M3_M2_CDNS_765593305589 $T=78120 186000 0 0 $X=78040 $Y=185870
X414 62 M3_M2_CDNS_765593305589 $T=78720 184820 0 0 $X=78640 $Y=184690
X415 104 M3_M2_CDNS_765593305589 $T=79890 191610 0 0 $X=79810 $Y=191480
X416 59 M3_M2_CDNS_765593305589 $T=80240 191340 0 0 $X=80160 $Y=191210
X417 31 M3_M2_CDNS_765593305589 $T=82410 190150 0 0 $X=82330 $Y=190020
X418 63 M3_M2_CDNS_765593305589 $T=82430 180700 0 0 $X=82350 $Y=180570
X419 91 M3_M2_CDNS_765593305589 $T=82800 188100 0 0 $X=82720 $Y=187970
X420 92 M3_M2_CDNS_765593305589 $T=83710 185900 0 0 $X=83630 $Y=185770
X421 65 M3_M2_CDNS_765593305589 $T=84170 177850 0 0 $X=84090 $Y=177720
X422 15 M3_M2_CDNS_765593305589 $T=84810 189220 0 0 $X=84730 $Y=189090
X423 40 M3_M2_CDNS_765593305589 $T=85640 186730 0 0 $X=85560 $Y=186600
X424 112 M3_M2_CDNS_765593305589 $T=91420 190110 0 0 $X=91340 $Y=189980
X425 42 M3_M2_CDNS_765593305589 $T=96230 190380 0 0 $X=96150 $Y=190250
X426 91 M3_M2_CDNS_765593305589 $T=96730 187430 0 0 $X=96650 $Y=187300
X427 89 M3_M2_CDNS_765593305589 $T=97030 190200 0 0 $X=96950 $Y=190070
X428 94 M4_M3_CDNS_7655933055810 $T=38650 183500 0 0 $X=38520 $Y=183420
X429 88 M4_M3_CDNS_7655933055810 $T=39000 187750 0 0 $X=38870 $Y=187670
X430 36 M4_M3_CDNS_7655933055810 $T=43110 170800 0 0 $X=42980 $Y=170720
X431 21 M4_M3_CDNS_7655933055810 $T=43950 190600 0 0 $X=43820 $Y=190520
X432 62 M4_M3_CDNS_7655933055810 $T=44650 184650 0 0 $X=44520 $Y=184570
X433 79 M4_M3_CDNS_7655933055810 $T=45000 185000 0 0 $X=44870 $Y=184920
X434 22 M4_M3_CDNS_7655933055810 $T=45350 185600 0 0 $X=45220 $Y=185520
X435 59 M4_M3_CDNS_7655933055810 $T=46050 185300 0 0 $X=45920 $Y=185220
X436 81 M4_M3_CDNS_7655933055810 $T=46400 183850 0 0 $X=46270 $Y=183770
X437 104 M4_M3_CDNS_7655933055810 $T=48860 182500 0 0 $X=48730 $Y=182420
X438 33 M4_M3_CDNS_7655933055810 $T=51340 188470 0 0 $X=51210 $Y=188390
X439 107 M4_M3_CDNS_7655933055810 $T=52210 183200 0 0 $X=52080 $Y=183120
X440 14 M4_M3_CDNS_7655933055810 $T=52840 161950 0 0 $X=52710 $Y=161870
X441 34 M4_M3_CDNS_7655933055810 $T=53210 175750 0 0 $X=53080 $Y=175670
X442 11 M4_M3_CDNS_7655933055810 $T=53630 182800 0 0 $X=53500 $Y=182720
X443 94 M4_M3_CDNS_7655933055810 $T=53630 183500 0 0 $X=53500 $Y=183420
X444 81 M4_M3_CDNS_7655933055810 $T=53630 183850 0 0 $X=53500 $Y=183770
X445 6 M4_M3_CDNS_7655933055810 $T=53630 184200 0 0 $X=53500 $Y=184120
X446 22 M4_M3_CDNS_7655933055810 $T=53630 185600 0 0 $X=53500 $Y=185520
X447 39 M4_M3_CDNS_7655933055810 $T=54830 189190 0 0 $X=54700 $Y=189110
X448 1 M4_M3_CDNS_7655933055810 $T=54990 178190 0 0 $X=54860 $Y=178110
X449 31 M4_M3_CDNS_7655933055810 $T=55250 189150 0 0 $X=55120 $Y=189070
X450 84 M4_M3_CDNS_7655933055810 $T=56210 188050 0 0 $X=56080 $Y=187970
X451 39 M4_M3_CDNS_7655933055810 $T=57000 170690 0 0 $X=56870 $Y=170610
X452 109 M4_M3_CDNS_7655933055810 $T=58750 188100 0 0 $X=58620 $Y=188020
X453 80 M4_M3_CDNS_7655933055810 $T=60980 186700 0 0 $X=60850 $Y=186620
X454 86 M4_M3_CDNS_7655933055810 $T=61520 199460 0 0 $X=61390 $Y=199380
X455 40 M4_M3_CDNS_7655933055810 $T=62060 186700 0 0 $X=61930 $Y=186620
X456 42 M4_M3_CDNS_7655933055810 $T=62230 187400 0 0 $X=62100 $Y=187320
X457 82 M4_M3_CDNS_7655933055810 $T=62320 202620 0 0 $X=62190 $Y=202540
X458 27 M4_M3_CDNS_7655933055810 $T=63360 190140 0 0 $X=63230 $Y=190060
X459 112 M4_M3_CDNS_7655933055810 $T=63730 190900 0 0 $X=63600 $Y=190820
X460 88 M4_M3_CDNS_7655933055810 $T=66160 187750 0 0 $X=66030 $Y=187670
X461 33 M4_M3_CDNS_7655933055810 $T=66830 182800 0 0 $X=66700 $Y=182720
X462 21 M4_M3_CDNS_7655933055810 $T=67650 190600 0 0 $X=67520 $Y=190520
X463 24 M4_M3_CDNS_7655933055810 $T=70970 169090 0 0 $X=70840 $Y=169010
X464 24 M4_M3_CDNS_7655933055810 $T=70970 190580 0 0 $X=70840 $Y=190500
X465 32 M4_M3_CDNS_7655933055810 $T=71630 189500 0 0 $X=71500 $Y=189420
X466 34 M4_M3_CDNS_7655933055810 $T=73630 175750 0 0 $X=73500 $Y=175670
X467 65 M4_M3_CDNS_7655933055810 $T=75630 175400 0 0 $X=75500 $Y=175320
X468 38 M4_M3_CDNS_7655933055810 $T=77010 183900 0 0 $X=76880 $Y=183820
X469 83 M4_M3_CDNS_7655933055810 $T=77510 185600 0 0 $X=77380 $Y=185520
X470 13 M4_M3_CDNS_7655933055810 $T=78460 190200 0 0 $X=78330 $Y=190120
X471 31 M4_M3_CDNS_7655933055810 $T=82410 189150 0 0 $X=82280 $Y=189070
X472 91 M4_M3_CDNS_7655933055810 $T=82800 189730 0 0 $X=82670 $Y=189650
X473 15 M4_M3_CDNS_7655933055810 $T=84810 188450 0 0 $X=84680 $Y=188370
X474 122 M3_M2_CDNS_7655933055811 $T=41130 153500 0 0 $X=41000 $Y=153370
X475 41 M3_M2_CDNS_7655933055811 $T=58340 152150 0 0 $X=58210 $Y=152020
X476 128 M3_M2_CDNS_7655933055811 $T=67780 149140 0 0 $X=67650 $Y=149010
X477 97 M3_M2_CDNS_7655933055811 $T=73560 153330 0 0 $X=73430 $Y=153200
X478 86 M3_M2_CDNS_7655933055812 $T=36550 200380 0 0 $X=36300 $Y=200300
X479 109 M3_M2_CDNS_7655933055812 $T=56450 200950 0 0 $X=56200 $Y=200870
X480 105 M3_M2_CDNS_7655933055812 $T=57700 162210 0 0 $X=57450 $Y=162130
X481 42 M3_M2_CDNS_7655933055812 $T=62230 187080 0 0 $X=61980 $Y=187000
X482 127 M3_M2_CDNS_7655933055812 $T=67160 148490 0 0 $X=66910 $Y=148410
X483 127 M3_M2_CDNS_7655933055813 $T=67370 152380 0 0 $X=67240 $Y=152250
X484 128 M3_M2_CDNS_7655933055813 $T=67820 152730 0 0 $X=67690 $Y=152600
X485 34 M4_M3_CDNS_7655933055814 $T=53210 177850 0 0 $X=53080 $Y=177720
X486 79 M4_M3_CDNS_7655933055814 $T=53420 186300 0 0 $X=53290 $Y=186170
X487 83 M4_M3_CDNS_7655933055814 $T=55950 186300 0 0 $X=55820 $Y=186170
X488 108 M4_M3_CDNS_7655933055814 $T=57350 169570 0 0 $X=57220 $Y=169440
X489 85 M4_M3_CDNS_7655933055814 $T=57590 186350 0 0 $X=57460 $Y=186220
X490 59 M4_M3_CDNS_7655933055814 $T=80240 191340 0 0 $X=80110 $Y=191210
X491 11 M4_M3_CDNS_7655933055815 $T=38220 182800 0 0 $X=38140 $Y=182670
X492 78 M4_M3_CDNS_7655933055815 $T=39970 182100 0 0 $X=39890 $Y=181970
X493 16 M4_M3_CDNS_7655933055815 $T=42200 171820 0 0 $X=42120 $Y=171690
X494 16 M4_M3_CDNS_7655933055815 $T=42200 176870 0 0 $X=42120 $Y=176740
X495 102 M4_M3_CDNS_7655933055815 $T=44700 185950 0 0 $X=44620 $Y=185820
X496 27 M4_M3_CDNS_7655933055815 $T=47120 190140 0 0 $X=47040 $Y=190010
X497 103 M4_M3_CDNS_7655933055815 $T=47510 163650 0 0 $X=47430 $Y=163520
X498 14 M4_M3_CDNS_7655933055815 $T=52840 180960 0 0 $X=52760 $Y=180830
X499 1 M4_M3_CDNS_7655933055815 $T=53500 189790 0 0 $X=53420 $Y=189660
X500 105 M4_M3_CDNS_7655933055815 $T=57700 162570 0 0 $X=57620 $Y=162440
X501 49 M4_M3_CDNS_7655933055815 $T=67710 190250 0 0 $X=67630 $Y=190120
X502 78 M4_M3_CDNS_7655933055815 $T=78120 182100 0 0 $X=78040 $Y=181970
X503 99 M4_M3_CDNS_7655933055815 $T=82040 188080 0 0 $X=81960 $Y=187950
X504 85 M4_M3_CDNS_7655933055815 $T=83580 186700 0 0 $X=83500 $Y=186570
X505 112 M4_M3_CDNS_7655933055815 $T=91420 190900 0 0 $X=91340 $Y=190770
X506 42 M4_M3_CDNS_7655933055815 $T=96230 190120 0 0 $X=96150 $Y=189990
X507 102 M3_M2_CDNS_7655933055816 $T=44700 186580 0 0 $X=44330 $Y=186450
X508 14 M3_M2_CDNS_7655933055816 $T=52630 161950 0 0 $X=52260 $Y=161820
X509 34 M3_M2_CDNS_7655933055816 $T=53210 177850 0 0 $X=52840 $Y=177720
X510 29 M3_M2_CDNS_7655933055816 $T=56870 161900 0 0 $X=56500 $Y=161770
X511 4 M3_M2_CDNS_7655933055816 $T=61490 162160 0 0 $X=61120 $Y=162030
X512 39 M3_M2_CDNS_7655933055816 $T=61490 169570 0 0 $X=61120 $Y=169440
X513 6 M4_M3_CDNS_7655933055817 $T=35930 184200 0 0 $X=35800 $Y=183830
X514 99 M4_M3_CDNS_7655933055817 $T=39350 187050 0 0 $X=39220 $Y=186680
X515 9 M4_M3_CDNS_7655933055817 $T=44630 161500 0 0 $X=44500 $Y=161130
X516 103 M4_M3_CDNS_7655933055817 $T=47510 178550 0 0 $X=47380 $Y=178180
X517 82 M4_M3_CDNS_7655933055817 $T=50150 201310 0 0 $X=50020 $Y=200940
X518 105 M4_M3_CDNS_7655933055817 $T=53150 207870 0 0 $X=53020 $Y=207500
X519 15 M4_M3_CDNS_7655933055817 $T=53630 188450 0 0 $X=53500 $Y=188080
X520 108 M4_M3_CDNS_7655933055817 $T=53890 207420 0 0 $X=53760 $Y=207050
X521 32 M4_M3_CDNS_7655933055817 $T=53900 189500 0 0 $X=53770 $Y=189130
X522 3 M4_M3_CDNS_7655933055817 $T=55250 191340 0 0 $X=55120 $Y=190970
X523 38 M4_M3_CDNS_7655933055817 $T=56450 192730 0 0 $X=56320 $Y=192360
X524 109 M4_M3_CDNS_7655933055817 $T=56450 200950 0 0 $X=56320 $Y=200580
X525 98 M4_M3_CDNS_7655933055817 $T=59010 188800 0 0 $X=58880 $Y=188430
X526 4 M4_M3_CDNS_7655933055817 $T=61490 162160 0 0 $X=61360 $Y=161790
X527 102 M4_M3_CDNS_7655933055817 $T=77510 189900 0 0 $X=77380 $Y=189530
X528 107 M4_M3_CDNS_7655933055817 $T=78220 189850 0 0 $X=78090 $Y=189480
X529 84 M4_M3_CDNS_7655933055817 $T=78690 189850 0 0 $X=78560 $Y=189480
X530 62 M4_M3_CDNS_7655933055817 $T=78720 184650 0 0 $X=78590 $Y=184280
X531 91 M4_M3_CDNS_7655933055817 $T=79550 189730 0 0 $X=79420 $Y=189360
X532 104 M4_M3_CDNS_7655933055817 $T=79890 191610 0 0 $X=79760 $Y=191240
X533 65 M4_M3_CDNS_7655933055817 $T=84170 177850 0 0 $X=84040 $Y=177480
X534 86 M4_M3_CDNS_7655933055818 $T=36550 200380 0 0 $X=36300 $Y=200300
X535 98 M4_M3_CDNS_7655933055818 $T=59010 172200 0 0 $X=58760 $Y=172120
X536 9 M4_M3_CDNS_7655933055818 $T=65000 181400 0 0 $X=64750 $Y=181320
X537 13 M4_M3_CDNS_7655933055818 $T=65630 179250 0 0 $X=65380 $Y=179170
X538 49 M4_M3_CDNS_7655933055818 $T=67710 172550 0 0 $X=67460 $Y=172470
X539 33 M5_M4_CDNS_7655933055820 $T=54050 184200 0 0 $X=53920 $Y=184120
X540 84 M5_M4_CDNS_7655933055820 $T=55600 183600 0 0 $X=55470 $Y=183520
X541 84 M5_M4_CDNS_7655933055820 $T=55600 188050 0 0 $X=55470 $Y=187970
X542 83 M5_M4_CDNS_7655933055820 $T=55950 185600 0 0 $X=55820 $Y=185520
X543 39 M5_M4_CDNS_7655933055820 $T=56300 170690 0 0 $X=56170 $Y=170610
X544 105 M5_M4_CDNS_7655933055820 $T=57700 179000 0 0 $X=57570 $Y=178920
X545 109 M5_M4_CDNS_7655933055820 $T=58050 200950 0 0 $X=57920 $Y=200870
X546 80 M5_M4_CDNS_7655933055820 $T=60980 180000 0 0 $X=60850 $Y=179920
X547 33 M5_M4_CDNS_7655933055820 $T=66830 184200 0 0 $X=66700 $Y=184120
X548 49 M5_M4_CDNS_7655933055820 $T=67710 189800 0 0 $X=67580 $Y=189720
X549 13 M5_M4_CDNS_7655933055820 $T=69630 190200 0 0 $X=69500 $Y=190120
X550 38 M5_M4_CDNS_7655933055820 $T=77010 192730 0 0 $X=76880 $Y=192650
X551 102 M5_M4_CDNS_7655933055820 $T=77510 185950 0 0 $X=77380 $Y=185870
X552 99 M5_M4_CDNS_7655933055820 $T=82040 187050 0 0 $X=81910 $Y=186970
X553 98 M5_M4_CDNS_7655933055821 $T=59010 172200 0 0 $X=58760 $Y=172120
X554 13 M5_M4_CDNS_7655933055821 $T=65630 179250 0 0 $X=65380 $Y=179170
X555 49 M5_M4_CDNS_7655933055821 $T=67710 172550 0 0 $X=67460 $Y=172470
X556 2 M5_M4_CDNS_7655933055822 $T=54550 200840 0 0 $X=54470 $Y=200590
X557 2 M5_M4_CDNS_7655933055822 $T=56650 178900 0 0 $X=56570 $Y=178650
X558 122 M2_M1_CDNS_7655933055823 $T=36060 146980 0 0 $X=35930 $Y=146850
X559 100 M2_M1_CDNS_7655933055823 $T=37190 148770 0 0 $X=37060 $Y=148640
X560 132 M2_M1_CDNS_7655933055823 $T=40240 148210 0 0 $X=40110 $Y=148080
X561 122 M2_M1_CDNS_7655933055823 $T=41060 147800 0 0 $X=40930 $Y=147670
X562 18 M2_M1_CDNS_7655933055823 $T=41550 210470 0 0 $X=41420 $Y=210340
X563 132 M2_M1_CDNS_7655933055823 $T=44780 154450 0 0 $X=44650 $Y=154320
X564 133 M2_M1_CDNS_7655933055823 $T=48770 148640 0 0 $X=48640 $Y=148510
X565 133 M2_M1_CDNS_7655933055823 $T=48770 154450 0 0 $X=48640 $Y=154320
X566 125 M2_M1_CDNS_7655933055823 $T=53670 149540 0 0 $X=53540 $Y=149410
X567 124 M2_M1_CDNS_7655933055823 $T=55200 149720 0 0 $X=55070 $Y=149590
X568 41 M2_M1_CDNS_7655933055823 $T=59140 149330 0 0 $X=59010 $Y=149200
X569 126 M2_M1_CDNS_7655933055823 $T=66860 154510 0 0 $X=66730 $Y=154380
X570 128 M2_M1_CDNS_7655933055823 $T=67820 153840 0 0 $X=67690 $Y=153710
X571 97 M2_M1_CDNS_7655933055823 $T=71450 149330 0 0 $X=71320 $Y=149200
X572 134 M2_M1_CDNS_7655933055823 $T=75890 149140 0 0 $X=75760 $Y=149010
X573 134 M2_M1_CDNS_7655933055823 $T=75890 154200 0 0 $X=75760 $Y=154070
X574 115 M2_M1_CDNS_7655933055823 $T=80260 149560 0 0 $X=80130 $Y=149430
X575 129 M2_M1_CDNS_7655933055823 $T=81770 149200 0 0 $X=81640 $Y=149070
X576 117 M2_M1_CDNS_7655933055823 $T=85850 149580 0 0 $X=85720 $Y=149450
X577 66 M2_M1_CDNS_7655933055823 $T=94350 149710 0 0 $X=94220 $Y=149580
X578 131 M2_M1_CDNS_7655933055823 $T=97100 142180 0 0 $X=96970 $Y=142050
X579 135 M2_M1_CDNS_7655933055823 $T=97460 141010 0 0 $X=97330 $Y=140880
X580 135 M2_M1_CDNS_7655933055823 $T=97460 154990 0 0 $X=97330 $Y=154860
X581 33 M5_M4_CDNS_7655933055824 $T=51340 188470 0 0 $X=51210 $Y=188100
X582 14 M5_M4_CDNS_7655933055824 $T=52840 180960 0 0 $X=52710 $Y=180590
X583 105 M5_M4_CDNS_7655933055824 $T=53150 207870 0 0 $X=53020 $Y=207500
X584 108 M5_M4_CDNS_7655933055824 $T=53890 207420 0 0 $X=53760 $Y=207050
X585 1 M5_M4_CDNS_7655933055824 $T=54990 178190 0 0 $X=54860 $Y=177820
X586 108 M5_M4_CDNS_7655933055824 $T=57350 169570 0 0 $X=57220 $Y=169200
X587 4 M5_M4_CDNS_7655933055824 $T=61490 162160 0 0 $X=61360 $Y=161790
X588 24 M5_M4_CDNS_7655933055824 $T=70970 169090 0 0 $X=70840 $Y=168720
X589 107 M5_M4_CDNS_7655933055824 $T=78220 189850 0 0 $X=78090 $Y=189480
X590 84 M5_M4_CDNS_7655933055824 $T=78690 189850 0 0 $X=78560 $Y=189480
X591 104 M5_M4_CDNS_7655933055824 $T=79890 191610 0 0 $X=79760 $Y=191240
X592 79 M5_M4_CDNS_7655933055825 $T=45000 186300 0 0 $X=44920 $Y=186170
X593 1 M5_M4_CDNS_7655933055825 $T=53500 189530 0 0 $X=53420 $Y=189400
X594 109 M5_M4_CDNS_7655933055825 $T=58050 188100 0 0 $X=57970 $Y=187970
X595 4 M5_M4_CDNS_7655933055825 $T=61490 209480 0 0 $X=61410 $Y=209350
X596 107 M5_M4_CDNS_7655933055825 $T=78220 183200 0 0 $X=78140 $Y=183070
X597 84 M5_M4_CDNS_7655933055825 $T=78690 183600 0 0 $X=78610 $Y=183470
X598 104 M5_M4_CDNS_7655933055825 $T=79890 182500 0 0 $X=79810 $Y=182370
X599 59 M5_M4_CDNS_7655933055825 $T=80240 185300 0 0 $X=80160 $Y=185170
X600 99 M5_M4_CDNS_7655933055825 $T=82040 187820 0 0 $X=81960 $Y=187690
X601 36 M4_M3_CDNS_7655933055828 $T=43110 179550 0 0 $X=42740 $Y=179420
X602 80 M4_M3_CDNS_7655933055828 $T=46270 179600 0 0 $X=45900 $Y=179470
X603 34 M4_M3_CDNS_7655933055828 $T=73630 178350 0 0 $X=73260 $Y=178220
X604 40 M4_M3_CDNS_7655933055828 $T=85640 186730 0 0 $X=85270 $Y=186600
X605 93 M2_M1_CDNS_7655933055829 $T=36870 154210 0 0 $X=36790 $Y=153960
X606 94 M2_M1_CDNS_7655933055829 $T=39090 200490 0 0 $X=39010 $Y=200240
X607 95 M2_M1_CDNS_7655933055829 $T=43880 210410 0 0 $X=43800 $Y=210160
X608 93 M2_M1_CDNS_7655933055829 $T=48210 153790 0 0 $X=48130 $Y=153540
X609 96 M2_M1_CDNS_7655933055829 $T=53980 160640 0 0 $X=53900 $Y=160390
X610 93 M2_M1_CDNS_7655933055829 $T=59550 153740 0 0 $X=59470 $Y=153490
X611 2 M2_M1_CDNS_7655933055829 $T=61490 178760 0 0 $X=61410 $Y=178510
X612 96 M2_M1_CDNS_7655933055829 $T=65090 160640 0 0 $X=65010 $Y=160390
X613 93 M2_M1_CDNS_7655933055829 $T=70770 153700 0 0 $X=70690 $Y=153450
X614 96 M2_M1_CDNS_7655933055829 $T=76650 169330 0 0 $X=76570 $Y=169080
X615 93 M2_M1_CDNS_7655933055829 $T=82230 153680 0 0 $X=82150 $Y=153430
X616 96 M2_M1_CDNS_7655933055829 $T=87810 169220 0 0 $X=87730 $Y=168970
X617 93 M2_M1_CDNS_7655933055829 $T=93570 153650 0 0 $X=93490 $Y=153400
X618 79 M5_M4_CDNS_7655933055830 $T=45000 185000 0 0 $X=44870 $Y=184870
X619 14 M5_M4_CDNS_7655933055830 $T=52840 161950 0 0 $X=52710 $Y=161820
X620 83 M5_M4_CDNS_7655933055830 $T=55950 186300 0 0 $X=55820 $Y=186170
X621 59 M5_M4_CDNS_7655933055830 $T=80240 191340 0 0 $X=80110 $Y=191210
X622 20 M3_M2_CDNS_7655933055831 $T=44740 169870 0 0 $X=44610 $Y=169740
X623 5 M3_M2_CDNS_7655933055831 $T=46030 163120 0 0 $X=45900 $Y=162990
X624 38 M3_M2_CDNS_7655933055831 $T=56450 192730 0 0 $X=56320 $Y=192600
X625 99 M3_M2_CDNS_7655933055831 $T=90620 191090 0 0 $X=90490 $Y=190960
X626 39 M5_M4_CDNS_7655933055832 $T=54830 189190 0 0 $X=54460 $Y=189060
X627 98 M5_M4_CDNS_7655933055832 $T=59010 188800 0 0 $X=58640 $Y=188670
X628 80 M5_M4_CDNS_7655933055832 $T=60980 186700 0 0 $X=60610 $Y=186570
X629 33 M5_M4_CDNS_7655933055832 $T=66830 182800 0 0 $X=66460 $Y=182670
X630 24 M5_M4_CDNS_7655933055832 $T=70970 190580 0 0 $X=70600 $Y=190450
X631 38 M5_M4_CDNS_7655933055832 $T=77010 183900 0 0 $X=76640 $Y=183770
X632 102 M5_M4_CDNS_7655933055832 $T=77510 189900 0 0 $X=77140 $Y=189770
X633 36 M3_M2_CDNS_7655933055833 $T=54580 170800 0 0 $X=54210 $Y=170720
X634 113 M3_M2_CDNS_7655933055833 $T=87620 190970 0 0 $X=87250 $Y=190890
X635 2 M4_M3_CDNS_7655933055836 $T=54550 200840 0 0 $X=54470 $Y=200590
X636 4 M3_M2_CDNS_7655933055838 $T=58900 209500 0 0 $X=58820 $Y=209250
X637 136 96 93 5 207 Diver $T=40660 207630 1 90 $X=36810 $Y=208360
X638 137 96 93 18 208 Diver $T=43640 207630 1 90 $X=39790 $Y=208360
X639 138 96 93 95 209 Diver $T=41440 207580 0 90 $X=42480 $Y=208310
X640 139 96 93 103 210 Diver $T=44420 207620 0 90 $X=45460 $Y=208350
X641 140 96 93 105 211 Diver $T=52000 207660 1 90 $X=48150 $Y=208390
X642 141 96 93 108 212 Diver $T=54980 207650 1 90 $X=51130 $Y=208380
X643 142 96 93 39 213 Diver $T=52780 207610 0 90 $X=53820 $Y=208340
X644 143 96 93 4 214 Diver $T=55760 207590 0 90 $X=56800 $Y=208320
X645 8 93 7 14 9 96 216 215 485 627
+ 628 486 HAdder $T=36010 162410 0 0 $X=36810 $Y=153450
X646 87 93 12 15 99 96 218 217 487 629
+ 630 488 HAdder $T=36010 188215 0 0 $X=36810 $Y=179255
X647 100 93 144 7 17 96 220 219 489 631
+ 632 490 HAdder $T=36010 194985 0 0 $X=36810 $Y=186025
X648 10 93 101 94 6 96 222 221 491 633
+ 634 492 HAdder $T=36010 201915 0 0 $X=36810 $Y=192955
X649 26 93 145 18 24 96 224 223 493 635
+ 636 494 HAdder $T=49070 171010 1 180 $X=42480 $Y=162050
X650 29 93 146 95 10 96 226 225 495 637
+ 638 496 HAdder $T=47350 171010 0 0 $X=48150 $Y=162050
X651 30 93 60 106 147 96 228 227 497 639
+ 640 498 HAdder $T=47350 179610 0 0 $X=48150 $Y=170650
X652 65 93 64 83 85 96 230 229 499 641
+ 642 500 HAdder $T=60410 188215 1 180 $X=53820 $Y=179255
X653 66 93 117 148 56 96 232 231 501 643
+ 644 502 HAdder $T=81370 162410 0 0 $X=82170 $Y=153450
X654 131 93 130 149 75 96 234 233 503 645
+ 646 504 HAdder $T=94430 162410 1 180 $X=87840 $Y=153450
X655 74 93 149 119 70 96 236 235 505 647
+ 648 506 HAdder $T=94430 171010 1 180 $X=87840 $Y=162050
X656 150 93 135 151 74 96 238 237 507 649
+ 650 508 HAdder $T=92710 162410 0 0 $X=93510 $Y=153450
X657 152 93 151 153 77 96 240 239 509 651
+ 652 510 HAdder $T=92710 171010 0 0 $X=93510 $Y=162050
X658 154 93 153 155 121 96 242 241 511 653
+ 654 512 HAdder $T=92710 179610 0 0 $X=93510 $Y=170650
X659 156 93 155 157 76 96 244 243 513 655
+ 656 514 HAdder $T=92710 188210 0 0 $X=93510 $Y=179250
X660 158 159 160 161 162 163 164 165 166 96
+ 93 89 91 68 73 157 167 168 42 50
+ 90 120 69 71 76 169 99 112 57 52
+ 113 61 116 72 170 63 15 40 13 62
+ 31 85 92 171 59 104 84 38 78 102
+ 107 83 172 6 22 32 28 111 88 27
+ 3 173 24 94 25 33 109 49 21 106
+ 174 9 11 79 81 82 110 98 80 17
+ 14 86 WallaceMultiplier $T=103430 160340 1 180 $X=59490 $Y=190900
X661 93 20 49 51 98 175 96 311 310 309 FAdder $T=35720 171510 1 0 $X=36810 $Y=162050
X662 93 16 78 175 88 13 96 314 313 312 FAdder $T=35720 180110 1 0 $X=36810 $Y=170650
X663 93 137 11 136 86 101 96 317 316 315 FAdder $T=35720 199385 0 0 $X=36810 $Y=200245
X664 93 122 145 132 5 8 96 320 319 318 FAdder $T=49360 162910 0 180 $X=42480 $Y=153450
X665 93 53 21 23 80 176 96 323 322 321 FAdder $T=49360 180110 0 180 $X=42480 $Y=170650
X666 93 19 102 176 27 62 96 326 325 324 FAdder $T=49360 188715 0 180 $X=42480 $Y=179255
X667 93 36 22 177 25 59 96 329 328 327 FAdder $T=49360 192095 1 180 $X=42480 $Y=192955
X668 93 138 79 139 81 177 96 332 331 330 FAdder $T=49360 199385 1 180 $X=42480 $Y=200245
X669 93 123 146 133 103 26 96 335 334 333 FAdder $T=47060 162910 1 0 $X=48150 $Y=153450
X670 93 34 107 147 3 31 96 338 337 336 FAdder $T=47060 188715 1 0 $X=48150 $Y=179255
X671 93 1 32 178 28 104 96 341 340 339 FAdder $T=47060 192095 0 0 $X=48150 $Y=192955
X672 93 141 33 140 82 178 96 344 343 342 FAdder $T=47060 199385 0 0 $X=48150 $Y=200245
X673 93 124 179 125 105 29 96 347 346 345 FAdder $T=60700 162910 0 180 $X=53820 $Y=153450
X674 93 35 180 179 108 36 96 350 349 348 FAdder $T=60700 171510 0 180 $X=53820 $Y=162050
X675 93 37 12 180 1 63 96 353 352 351 FAdder $T=60700 180110 0 180 $X=53820 $Y=170650
X676 93 2 38 181 111 84 96 356 355 354 FAdder $T=60700 192095 1 180 $X=53820 $Y=192955
X677 93 142 109 143 110 181 96 359 358 357 FAdder $T=60700 199385 1 180 $X=53820 $Y=200245
X678 93 127 182 41 4 35 96 362 361 360 FAdder $T=58400 162910 1 0 $X=59490 $Y=153450
X679 93 43 183 182 39 37 96 365 364 363 FAdder $T=58400 171510 1 0 $X=59490 $Y=162050
X680 93 44 184 183 2 87 96 368 367 366 FAdder $T=58400 180110 1 0 $X=59490 $Y=170650
X681 93 45 112 184 40 42 96 371 370 369 FAdder $T=58400 188715 1 0 $X=59490 $Y=179255
X682 93 128 185 126 51 43 96 374 373 372 FAdder $T=72040 162910 0 180 $X=65160 $Y=153450
X683 93 46 186 185 20 44 96 377 376 375 FAdder $T=72040 171510 0 180 $X=65160 $Y=162050
X684 93 47 187 186 16 45 96 380 379 378 FAdder $T=72040 180110 0 180 $X=65160 $Y=170650
X685 93 48 57 187 52 50 96 383 382 381 FAdder $T=72040 188715 0 180 $X=65160 $Y=179255
X686 93 134 188 97 23 46 96 386 385 384 FAdder $T=69740 162910 1 0 $X=70830 $Y=153450
X687 93 54 189 188 53 47 96 389 388 387 FAdder $T=69740 171510 1 0 $X=70830 $Y=162050
X688 93 55 190 189 19 48 96 392 391 390 FAdder $T=69740 180110 1 0 $X=70830 $Y=170650
X689 93 58 90 190 113 89 96 395 394 393 FAdder $T=69740 188715 1 0 $X=70830 $Y=179255
X690 93 129 191 115 60 54 96 398 397 396 FAdder $T=83380 162910 0 180 $X=76500 $Y=153450
X691 93 56 192 191 30 55 96 401 400 399 FAdder $T=83380 171510 0 180 $X=76500 $Y=162050
X692 93 114 193 192 34 58 96 404 403 402 FAdder $T=83380 180110 0 180 $X=76500 $Y=170650
X693 93 67 120 193 61 91 96 407 406 405 FAdder $T=83380 188715 0 180 $X=76500 $Y=179255
X694 93 75 194 148 64 114 96 410 409 408 FAdder $T=81080 171510 1 0 $X=82170 $Y=162050
X695 93 70 195 194 65 67 96 413 412 411 FAdder $T=81080 180110 1 0 $X=82170 $Y=170650
X696 93 118 69 195 116 68 96 416 415 414 FAdder $T=81080 188715 1 0 $X=82170 $Y=179255
X697 93 77 196 119 92 118 96 419 418 417 FAdder $T=94720 180110 0 180 $X=87840 $Y=170650
X698 93 121 71 196 72 73 96 422 421 420 FAdder $T=94720 188710 0 180 $X=87840 $Y=179250
X699 122 132 100 197 93 96 133 198 123 125
+ 199 124 41 200 126 201 127 128 97 202
+ 134 115 203 129 117 204 205 130 206 66
+ 131 135 423 440 444 449 432 468 472 477
+ 426 434 438 436 433 462 466 464 461 460
+ 425 427 430 431 455 457 458 459 WallaceFinalAdder $T=36320 132010 0 0 $X=36320 $Y=132010
M0 207 136 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=37590 $Y=208970 $dt=0
M1 5 207 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=37590 $Y=209900 $dt=0
M2 51 309 49 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=163470 $dt=0
M3 20 309 175 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=164810 $dt=0
M4 309 175 20 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=165220 $dt=0
M5 311 49 310 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=166150 $dt=0
M6 49 310 311 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=166560 $dt=0
M7 309 98 49 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=166970 $dt=0
M8 98 49 309 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=167380 $dt=0
M9 175 312 78 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=172070 $dt=0
M10 16 312 13 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=173410 $dt=0
M11 312 13 16 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=173820 $dt=0
M12 314 78 313 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=174750 $dt=0
M13 78 313 314 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=175160 $dt=0
M14 312 88 78 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=175570 $dt=0
M15 88 78 312 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=175980 $dt=0
M16 315 11 86 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=203425 $dt=0
M17 11 86 315 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=203835 $dt=0
M18 317 316 11 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=204245 $dt=0
M19 316 11 317 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=204655 $dt=0
M20 137 101 315 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=205585 $dt=0
M21 101 315 137 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=205995 $dt=0
M22 11 315 136 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=37700 $Y=207335 $dt=0
M23 208 137 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=40570 $Y=208970 $dt=0
M24 18 208 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=40570 $Y=209900 $dt=0
M25 209 138 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=44270 $Y=208920 $dt=0
M26 95 209 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=44270 $Y=209850 $dt=0
M27 132 318 145 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=154870 $dt=0
M28 122 318 8 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=156210 $dt=0
M29 318 8 122 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=156620 $dt=0
M30 320 145 319 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=157550 $dt=0
M31 145 319 320 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=157960 $dt=0
M32 318 5 145 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=158370 $dt=0
M33 5 145 318 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=158780 $dt=0
M34 23 321 21 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=172070 $dt=0
M35 53 321 176 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=173410 $dt=0
M36 321 176 53 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=173820 $dt=0
M37 323 21 322 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=174750 $dt=0
M38 21 322 323 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=175160 $dt=0
M39 321 80 21 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=175570 $dt=0
M40 80 21 321 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=175980 $dt=0
M41 176 324 102 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=180675 $dt=0
M42 19 324 62 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=182015 $dt=0
M43 324 62 19 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=182425 $dt=0
M44 326 102 325 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=183355 $dt=0
M45 102 325 326 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=183765 $dt=0
M46 324 27 102 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=184175 $dt=0
M47 27 102 324 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=184585 $dt=0
M48 327 22 25 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=196135 $dt=0
M49 22 25 327 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=196545 $dt=0
M50 329 328 22 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=196955 $dt=0
M51 328 22 329 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=197365 $dt=0
M52 36 59 327 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=198295 $dt=0
M53 59 327 36 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=198705 $dt=0
M54 22 327 177 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=200045 $dt=0
M55 330 79 81 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=203425 $dt=0
M56 79 81 330 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=203835 $dt=0
M57 332 331 79 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=204245 $dt=0
M58 331 79 332 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=204655 $dt=0
M59 138 177 330 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=205585 $dt=0
M60 177 330 138 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=205995 $dt=0
M61 79 330 139 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=47140 $Y=207335 $dt=0
M62 210 139 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=47250 $Y=208960 $dt=0
M63 103 210 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=47250 $Y=209890 $dt=0
M64 211 140 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=48930 $Y=209000 $dt=0
M65 105 211 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=48930 $Y=209930 $dt=0
M66 133 333 146 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=154870 $dt=0
M67 123 333 26 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=156210 $dt=0
M68 333 26 123 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=156620 $dt=0
M69 335 146 334 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=157550 $dt=0
M70 146 334 335 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=157960 $dt=0
M71 333 103 146 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=158370 $dt=0
M72 103 146 333 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=158780 $dt=0
M73 147 336 107 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=180675 $dt=0
M74 34 336 31 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=182015 $dt=0
M75 336 31 34 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=182425 $dt=0
M76 338 107 337 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=183355 $dt=0
M77 107 337 338 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=183765 $dt=0
M78 336 3 107 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=184175 $dt=0
M79 3 107 336 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=184585 $dt=0
M80 339 32 28 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=196135 $dt=0
M81 32 28 339 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=196545 $dt=0
M82 341 340 32 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=196955 $dt=0
M83 340 32 341 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=197365 $dt=0
M84 1 104 339 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=198295 $dt=0
M85 104 339 1 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=198705 $dt=0
M86 32 339 178 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=200045 $dt=0
M87 342 33 82 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=203425 $dt=0
M88 33 82 342 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=203835 $dt=0
M89 344 343 33 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=204245 $dt=0
M90 343 33 344 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=204655 $dt=0
M91 141 178 342 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=205585 $dt=0
M92 178 342 141 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=205995 $dt=0
M93 33 342 140 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=49040 $Y=207335 $dt=0
M94 212 141 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=51910 $Y=208990 $dt=0
M95 108 212 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=51910 $Y=209920 $dt=0
M96 213 142 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=55610 $Y=208950 $dt=0
M97 39 213 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=55610 $Y=209880 $dt=0
M98 125 345 179 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.10357 scb=0.000255666 scc=3.44804e-08 $X=58480 $Y=154870 $dt=0
M99 124 345 29 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=156210 $dt=0
M100 345 29 124 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=156620 $dt=0
M101 347 179 346 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=157550 $dt=0
M102 179 346 347 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=157960 $dt=0
M103 345 105 179 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=158370 $dt=0
M104 105 179 345 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=158780 $dt=0
M105 179 348 180 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=163470 $dt=0
M106 35 348 36 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=164810 $dt=0
M107 348 36 35 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=165220 $dt=0
M108 350 180 349 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=166150 $dt=0
M109 180 349 350 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=166560 $dt=0
M110 348 108 180 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=166970 $dt=0
M111 108 180 348 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=167380 $dt=0
M112 180 351 12 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=172070 $dt=0
M113 37 351 63 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=173410 $dt=0
M114 351 63 37 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=173820 $dt=0
M115 353 12 352 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=174750 $dt=0
M116 12 352 353 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=175160 $dt=0
M117 351 1 12 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=175570 $dt=0
M118 1 12 351 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=175980 $dt=0
M119 354 38 111 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=58480 $Y=196135 $dt=0
M120 38 111 354 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=58480 $Y=196545 $dt=0
M121 356 355 38 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=58480 $Y=196955 $dt=0
M122 355 38 356 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=197365 $dt=0
M123 2 84 354 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=198295 $dt=0
M124 84 354 2 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=198705 $dt=0
M125 38 354 181 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=200045 $dt=0
M126 357 109 110 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=203425 $dt=0
M127 109 110 357 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=203835 $dt=0
M128 359 358 109 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=204245 $dt=0
M129 358 109 359 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=4.11282 scb=0.000306462 scc=1.0989e-07 $X=58480 $Y=204655 $dt=0
M130 142 181 357 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=58480 $Y=205585 $dt=0
M131 181 357 142 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=58480 $Y=205995 $dt=0
M132 109 357 143 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=58480 $Y=207335 $dt=0
M133 214 143 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=58590 $Y=208930 $dt=0
M134 4 214 93 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8263 scb=0.00911451 scc=0.000207374 $X=58590 $Y=209860 $dt=0
M135 41 360 182 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=154870 $dt=0
M136 127 360 35 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=156210 $dt=0
M137 360 35 127 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=156620 $dt=0
M138 362 182 361 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=157550 $dt=0
M139 182 361 362 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=157960 $dt=0
M140 360 4 182 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=158370 $dt=0
M141 4 182 360 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=158780 $dt=0
M142 182 363 183 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=163470 $dt=0
M143 43 363 37 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=164810 $dt=0
M144 363 37 43 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=165220 $dt=0
M145 365 183 364 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=166150 $dt=0
M146 183 364 365 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=166560 $dt=0
M147 363 39 183 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=166970 $dt=0
M148 39 183 363 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=167380 $dt=0
M149 183 366 184 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=172070 $dt=0
M150 44 366 87 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=173410 $dt=0
M151 366 87 44 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=173820 $dt=0
M152 368 184 367 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=174750 $dt=0
M153 184 367 368 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=175160 $dt=0
M154 366 2 184 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=175570 $dt=0
M155 2 184 366 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=175980 $dt=0
M156 184 369 112 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=180675 $dt=0
M157 45 369 42 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=182015 $dt=0
M158 369 42 45 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=182425 $dt=0
M159 371 112 370 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=183355 $dt=0
M160 112 370 371 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=183765 $dt=0
M161 369 40 112 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=184175 $dt=0
M162 40 112 369 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=60380 $Y=184585 $dt=0
M163 126 372 185 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.10624 scb=0.000256891 scc=3.49982e-08 $X=69820 $Y=154870 $dt=0
M164 128 372 43 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=156210 $dt=0
M165 372 43 128 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=156620 $dt=0
M166 374 185 373 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=157550 $dt=0
M167 185 373 374 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=157960 $dt=0
M168 372 51 185 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=158370 $dt=0
M169 51 185 372 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=158780 $dt=0
M170 185 375 186 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=163470 $dt=0
M171 46 375 44 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=164810 $dt=0
M172 375 44 46 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=165220 $dt=0
M173 377 186 376 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=166150 $dt=0
M174 186 376 377 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=166560 $dt=0
M175 375 20 186 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=166970 $dt=0
M176 20 186 375 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=167380 $dt=0
M177 186 378 187 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=172070 $dt=0
M178 47 378 45 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=173410 $dt=0
M179 378 45 47 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=173820 $dt=0
M180 380 187 379 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=174750 $dt=0
M181 187 379 380 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=175160 $dt=0
M182 378 16 187 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=175570 $dt=0
M183 16 187 378 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=175980 $dt=0
M184 187 381 57 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=180675 $dt=0
M185 48 381 50 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=182015 $dt=0
M186 381 50 48 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=182425 $dt=0
M187 383 57 382 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=183355 $dt=0
M188 57 382 383 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=183765 $dt=0
M189 381 52 57 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=184175 $dt=0
M190 52 57 381 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=69820 $Y=184585 $dt=0
M191 97 384 188 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.71642 scb=0.000135303 scc=5.64513e-09 $X=71720 $Y=154870 $dt=0
M192 134 384 46 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=156210 $dt=0
M193 384 46 134 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=156620 $dt=0
M194 386 188 385 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=157550 $dt=0
M195 188 385 386 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=157960 $dt=0
M196 384 23 188 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=158370 $dt=0
M197 23 188 384 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=158780 $dt=0
M198 188 387 189 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=163470 $dt=0
M199 54 387 47 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=164810 $dt=0
M200 387 47 54 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=165220 $dt=0
M201 389 189 388 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=166150 $dt=0
M202 189 388 389 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=166560 $dt=0
M203 387 53 189 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=166970 $dt=0
M204 53 189 387 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=167380 $dt=0
M205 189 390 190 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=172070 $dt=0
M206 55 390 48 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=173410 $dt=0
M207 390 48 55 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=173820 $dt=0
M208 392 190 391 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=174750 $dt=0
M209 190 391 392 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=175160 $dt=0
M210 390 19 190 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=175570 $dt=0
M211 19 190 390 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=175980 $dt=0
M212 190 393 90 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=180675 $dt=0
M213 58 393 89 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=182015 $dt=0
M214 393 89 58 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=182425 $dt=0
M215 395 90 394 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=183355 $dt=0
M216 90 394 395 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=183765 $dt=0
M217 393 113 90 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=184175 $dt=0
M218 113 90 393 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=71720 $Y=184585 $dt=0
M219 115 396 191 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=154870 $dt=0
M220 129 396 54 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=156210 $dt=0
M221 396 54 129 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=156620 $dt=0
M222 398 191 397 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=157550 $dt=0
M223 191 397 398 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=157960 $dt=0
M224 396 60 191 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=158370 $dt=0
M225 60 191 396 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=158780 $dt=0
M226 191 399 192 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=163470 $dt=0
M227 56 399 55 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=164810 $dt=0
M228 399 55 56 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=165220 $dt=0
M229 401 192 400 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=166150 $dt=0
M230 192 400 401 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=166560 $dt=0
M231 399 30 192 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=166970 $dt=0
M232 30 192 399 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=167380 $dt=0
M233 192 402 193 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=172070 $dt=0
M234 114 402 58 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=173410 $dt=0
M235 402 58 114 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=173820 $dt=0
M236 404 193 403 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=174750 $dt=0
M237 193 403 404 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=175160 $dt=0
M238 402 34 193 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=175570 $dt=0
M239 34 193 402 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=175980 $dt=0
M240 193 405 120 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=180675 $dt=0
M241 67 405 91 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=182015 $dt=0
M242 405 91 67 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=182425 $dt=0
M243 407 120 406 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=183355 $dt=0
M244 120 406 407 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=183765 $dt=0
M245 405 61 120 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=184175 $dt=0
M246 61 120 405 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=81160 $Y=184585 $dt=0
M247 148 408 194 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=163470 $dt=0
M248 75 408 114 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=164810 $dt=0
M249 408 114 75 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=165220 $dt=0
M250 410 194 409 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=166150 $dt=0
M251 194 409 410 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=166560 $dt=0
M252 408 64 194 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=166970 $dt=0
M253 64 194 408 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=167380 $dt=0
M254 194 411 195 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=172070 $dt=0
M255 70 411 67 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=173410 $dt=0
M256 411 67 70 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=173820 $dt=0
M257 413 195 412 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=174750 $dt=0
M258 195 412 413 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=175160 $dt=0
M259 411 65 195 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=175570 $dt=0
M260 65 195 411 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=175980 $dt=0
M261 195 414 69 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=180675 $dt=0
M262 118 414 68 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=182015 $dt=0
M263 414 68 118 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=182425 $dt=0
M264 416 69 415 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=183355 $dt=0
M265 69 415 416 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=183765 $dt=0
M266 414 116 69 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=184175 $dt=0
M267 116 69 414 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=83060 $Y=184585 $dt=0
M268 119 417 196 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=172070 $dt=0
M269 77 417 118 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=173410 $dt=0
M270 417 118 77 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=173820 $dt=0
M271 419 196 418 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=174750 $dt=0
M272 196 418 419 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=175160 $dt=0
M273 417 92 196 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=175570 $dt=0
M274 92 196 417 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=175980 $dt=0
M275 196 420 71 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=180670 $dt=0
M276 121 420 73 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=182010 $dt=0
M277 420 73 121 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=182420 $dt=0
M278 422 71 421 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=183350 $dt=0
M279 71 421 422 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=183760 $dt=0
M280 420 72 71 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=184170 $dt=0
M281 72 71 420 93 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=92500 $Y=184580 $dt=0
M282 207 136 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=38600 $Y=208970 $dt=1
M283 5 207 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=38600 $Y=209900 $dt=1
M284 51 309 175 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=41150 $Y=163470 $dt=1
M285 175 312 13 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41150 $Y=172070 $dt=1
M286 101 315 136 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41150 $Y=207335 $dt=1
M287 628 216 7 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=41530 $Y=155520 $dt=1
M288 96 215 628 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=41530 $Y=155730 $dt=1
M289 96 215 627 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=41530 $Y=156660 $dt=1
M290 627 216 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=41530 $Y=157070 $dt=1
M291 8 9 627 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41530 $Y=157480 $dt=1
M292 627 14 8 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41530 $Y=157890 $dt=1
M293 96 14 215 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=41530 $Y=158820 $dt=1
M294 96 9 216 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=41530 $Y=159750 $dt=1
M295 630 218 12 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=41530 $Y=181325 $dt=1
M296 96 217 630 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=41530 $Y=181535 $dt=1
M297 96 217 629 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=41530 $Y=182465 $dt=1
M298 629 218 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=41530 $Y=182875 $dt=1
M299 87 99 629 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41530 $Y=183285 $dt=1
M300 629 15 87 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41530 $Y=183695 $dt=1
M301 96 15 217 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=41530 $Y=184625 $dt=1
M302 96 99 218 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=41530 $Y=185555 $dt=1
M303 632 220 144 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=41530 $Y=188095 $dt=1
M304 96 219 632 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=41530 $Y=188305 $dt=1
M305 96 219 631 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=41530 $Y=189235 $dt=1
M306 631 220 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=41530 $Y=189645 $dt=1
M307 100 17 631 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=41530 $Y=190055 $dt=1
M308 631 7 100 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=41530 $Y=190465 $dt=1
M309 96 7 219 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=41530 $Y=191395 $dt=1
M310 96 17 220 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=41530 $Y=192325 $dt=1
M311 634 222 101 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=41530 $Y=195025 $dt=1
M312 96 221 634 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=41530 $Y=195235 $dt=1
M313 96 221 633 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=41530 $Y=196165 $dt=1
M314 633 222 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=41530 $Y=196575 $dt=1
M315 10 6 633 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41530 $Y=196985 $dt=1
M316 633 94 10 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41530 $Y=197395 $dt=1
M317 96 94 221 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=41530 $Y=198325 $dt=1
M318 96 6 222 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=41530 $Y=199255 $dt=1
M319 208 137 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=41580 $Y=208970 $dt=1
M320 18 208 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=41580 $Y=209900 $dt=1
M321 209 138 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=43260 $Y=208920 $dt=1
M322 95 209 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=43260 $Y=209850 $dt=1
M323 636 224 145 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=43310 $Y=164120 $dt=1
M324 96 223 636 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=43310 $Y=164330 $dt=1
M325 96 223 635 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=43310 $Y=165260 $dt=1
M326 635 224 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=43310 $Y=165670 $dt=1
M327 26 24 635 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43310 $Y=166080 $dt=1
M328 635 18 26 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43310 $Y=166490 $dt=1
M329 96 18 223 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=43310 $Y=167420 $dt=1
M330 96 24 224 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=43310 $Y=168350 $dt=1
M331 132 318 8 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=43690 $Y=154870 $dt=1
M332 23 321 176 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=43690 $Y=172070 $dt=1
M333 176 324 62 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=43690 $Y=180675 $dt=1
M334 59 327 177 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=43690 $Y=200045 $dt=1
M335 177 330 139 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=43690 $Y=207335 $dt=1
M336 210 139 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=46240 $Y=208960 $dt=1
M337 103 210 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=46240 $Y=209890 $dt=1
M338 211 140 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=49940 $Y=209000 $dt=1
M339 105 211 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=49940 $Y=209930 $dt=1
M340 133 333 26 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52490 $Y=154870 $dt=1
M341 147 336 31 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=52490 $Y=180675 $dt=1
M342 104 339 178 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52490 $Y=200045 $dt=1
M343 178 342 140 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52490 $Y=207335 $dt=1
M344 638 226 146 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52870 $Y=164120 $dt=1
M345 96 225 638 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=52870 $Y=164330 $dt=1
M346 96 225 637 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=52870 $Y=165260 $dt=1
M347 637 226 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=52870 $Y=165670 $dt=1
M348 29 10 637 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52870 $Y=166080 $dt=1
M349 637 95 29 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52870 $Y=166490 $dt=1
M350 96 95 225 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=52870 $Y=167420 $dt=1
M351 96 10 226 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52870 $Y=168350 $dt=1
M352 640 228 60 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52870 $Y=172720 $dt=1
M353 96 227 640 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=52870 $Y=172930 $dt=1
M354 96 227 639 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=52870 $Y=173860 $dt=1
M355 639 228 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=52870 $Y=174270 $dt=1
M356 30 147 639 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52870 $Y=174680 $dt=1
M357 639 106 30 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52870 $Y=175090 $dt=1
M358 96 106 227 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=52870 $Y=176020 $dt=1
M359 96 147 228 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52870 $Y=176950 $dt=1
M360 212 141 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=52920 $Y=208990 $dt=1
M361 108 212 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=52920 $Y=209920 $dt=1
M362 213 142 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=54600 $Y=208950 $dt=1
M363 39 213 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=54600 $Y=209880 $dt=1
M364 642 230 64 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=54650 $Y=181325 $dt=1
M365 96 229 642 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=54650 $Y=181535 $dt=1
M366 96 229 641 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=54650 $Y=182465 $dt=1
M367 641 230 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=54650 $Y=182875 $dt=1
M368 65 85 641 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54650 $Y=183285 $dt=1
M369 641 83 65 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54650 $Y=183695 $dt=1
M370 96 83 229 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=54650 $Y=184625 $dt=1
M371 96 85 230 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=54650 $Y=185555 $dt=1
M372 125 345 29 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=55030 $Y=154870 $dt=1
M373 179 348 36 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=55030 $Y=163470 $dt=1
M374 180 351 63 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=55030 $Y=172070 $dt=1
M375 84 354 181 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=55030 $Y=200045 $dt=1
M376 181 357 143 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=55030 $Y=207335 $dt=1
M377 214 143 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=57580 $Y=208930 $dt=1
M378 4 214 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=57580 $Y=209860 $dt=1
M379 41 360 35 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=63830 $Y=154870 $dt=1
M380 182 363 37 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=63830 $Y=163470 $dt=1
M381 183 366 87 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=63830 $Y=172070 $dt=1
M382 184 369 42 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=63830 $Y=180675 $dt=1
M383 126 372 43 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=66370 $Y=154870 $dt=1
M384 185 375 44 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=66370 $Y=163470 $dt=1
M385 186 378 45 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=66370 $Y=172070 $dt=1
M386 187 381 50 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=66370 $Y=180675 $dt=1
M387 97 384 46 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=75170 $Y=154870 $dt=1
M388 188 387 47 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=75170 $Y=163470 $dt=1
M389 189 390 48 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=75170 $Y=172070 $dt=1
M390 190 393 89 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=75170 $Y=180675 $dt=1
M391 115 396 54 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=77710 $Y=154870 $dt=1
M392 191 399 55 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=77710 $Y=163470 $dt=1
M393 192 402 58 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=77710 $Y=172070 $dt=1
M394 193 405 91 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=77710 $Y=180675 $dt=1
M395 148 408 114 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=86510 $Y=163470 $dt=1
M396 194 411 67 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=86510 $Y=172070 $dt=1
M397 195 414 68 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=86510 $Y=180675 $dt=1
M398 644 232 117 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=86890 $Y=155520 $dt=1
M399 96 231 644 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.901 scb=0.0471116 scc=0.0116656 $X=86890 $Y=155730 $dt=1
M400 96 231 643 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.1268 scb=0.0349743 scc=0.0111863 $X=86890 $Y=156660 $dt=1
M401 643 232 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.5388 scb=0.0347327 scc=0.0111862 $X=86890 $Y=157070 $dt=1
M402 66 56 643 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=86890 $Y=157480 $dt=1
M403 643 148 66 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=86890 $Y=157890 $dt=1
M404 96 148 231 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.6513 scb=0.0354006 scc=0.011187 $X=86890 $Y=158820 $dt=1
M405 96 56 232 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=86890 $Y=159750 $dt=1
M406 646 234 130 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=88670 $Y=155520 $dt=1
M407 96 233 646 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.901 scb=0.0471116 scc=0.0116656 $X=88670 $Y=155730 $dt=1
M408 96 233 645 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.1268 scb=0.0349743 scc=0.0111863 $X=88670 $Y=156660 $dt=1
M409 645 234 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.5388 scb=0.0347327 scc=0.0111862 $X=88670 $Y=157070 $dt=1
M410 131 75 645 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=88670 $Y=157480 $dt=1
M411 645 149 131 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=88670 $Y=157890 $dt=1
M412 96 149 233 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.6513 scb=0.0354006 scc=0.011187 $X=88670 $Y=158820 $dt=1
M413 96 75 234 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=88670 $Y=159750 $dt=1
M414 648 236 149 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=88670 $Y=164120 $dt=1
M415 96 235 648 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=88670 $Y=164330 $dt=1
M416 96 235 647 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=88670 $Y=165260 $dt=1
M417 647 236 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=88670 $Y=165670 $dt=1
M418 74 70 647 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=88670 $Y=166080 $dt=1
M419 647 119 74 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=88670 $Y=166490 $dt=1
M420 96 119 235 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=88670 $Y=167420 $dt=1
M421 96 70 236 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=88670 $Y=168350 $dt=1
M422 119 417 118 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=89050 $Y=172070 $dt=1
M423 196 420 73 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=89050 $Y=180670 $dt=1
M424 650 238 135 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=155520 $dt=1
M425 96 237 650 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=98230 $Y=155730 $dt=1
M426 96 237 649 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=98230 $Y=156660 $dt=1
M427 649 238 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=98230 $Y=157070 $dt=1
M428 150 74 649 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=157480 $dt=1
M429 649 151 150 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=157890 $dt=1
M430 96 151 237 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=98230 $Y=158820 $dt=1
M431 96 74 238 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=159750 $dt=1
M432 652 240 151 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=164120 $dt=1
M433 96 239 652 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=98230 $Y=164330 $dt=1
M434 96 239 651 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=98230 $Y=165260 $dt=1
M435 651 240 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=98230 $Y=165670 $dt=1
M436 152 77 651 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=166080 $dt=1
M437 651 153 152 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=166490 $dt=1
M438 96 153 239 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=98230 $Y=167420 $dt=1
M439 96 77 240 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=168350 $dt=1
M440 654 242 153 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=172720 $dt=1
M441 96 241 654 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=98230 $Y=172930 $dt=1
M442 96 241 653 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=98230 $Y=173860 $dt=1
M443 653 242 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=98230 $Y=174270 $dt=1
M444 154 121 653 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=174680 $dt=1
M445 653 155 154 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=175090 $dt=1
M446 96 155 241 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=98230 $Y=176020 $dt=1
M447 96 121 242 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=176950 $dt=1
M448 656 244 155 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=181320 $dt=1
M449 96 243 656 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=98230 $Y=181530 $dt=1
M450 96 243 655 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=98230 $Y=182460 $dt=1
M451 655 244 96 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=98230 $Y=182870 $dt=1
M452 156 76 655 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=183280 $dt=1
M453 655 157 156 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=98230 $Y=183690 $dt=1
M454 96 157 243 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=98230 $Y=184620 $dt=1
M455 96 76 244 96 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=98230 $Y=185550 $dt=1
.ends WallaceProject
