* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : NAND                                         *
* Netlisted  : Mon Sep 22 20:30:35 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_758587431050                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_758587431050 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_758587431050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_758587431050                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_758587431050 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=125.222 scb=0.0727692 scc=0.0141076 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_758587431050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_758587431051                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_758587431051 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=5.13215 scb=0.00119239 scc=2.71899e-06 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_758587431051

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_758587431052                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_758587431052 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=125.222 scb=0.0727692 scc=0.0141076 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_758587431052

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_758587431053                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_758587431053 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=5.13215 scb=0.00119239 scc=2.71899e-06 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_758587431053

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND 5 1 2 4 3
** N=6 EP=5 FDC=4
X0 1 M1_PO_CDNS_758587431050 $T=580 -2090 0 90 $X=460 $Y=-2190
X1 2 M1_PO_CDNS_758587431050 $T=1460 -2100 0 90 $X=1340 $Y=-2200
X2 3 4 1 5 pmos1v_CDNS_758587431050 $T=840 -1460 0 0 $X=420 $Y=-1660
X3 5 2 6 nmos1v_CDNS_758587431051 $T=1340 -3130 1 180 $X=1050 $Y=-3970
X4 4 2 3 5 pmos1v_CDNS_758587431052 $T=1340 -1460 1 180 $X=1010 $Y=-1660
X5 3 1 6 5 nmos1v_CDNS_758587431053 $T=1130 -3130 1 180 $X=620 $Y=-3330
.ends NAND
