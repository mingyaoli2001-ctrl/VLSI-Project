* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 4bit_CLA_logic                               *
* Netlisted  : Sun Dec  7 11:09:58 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765123794260                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765123794260 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765123794260

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_765123794261                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_765123794261 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_765123794261

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765123794262                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765123794262 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765123794262

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765123794263                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765123794263 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765123794263

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765123794264                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765123794264 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765123794264

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_765123794265                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_765123794265 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_765123794265

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765123794266                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765123794266 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765123794266

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765123794267                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765123794267 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765123794267

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765123794268                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765123794268 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765123794268

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765123794269                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765123794269 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765123794269

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651237942610                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651237942610 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651237942610

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651237942611                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651237942611 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651237942611

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7651237942614                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7651237942614 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7651237942614

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651237942615                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651237942615 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651237942615

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7651237942616                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7651237942616 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7651237942616

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651237942617                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651237942617 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651237942617

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7651237942618                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7651237942618 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7651237942618

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7651237942619                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7651237942619 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7651237942619

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7651237942620                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7651237942620 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7651237942620

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7651237942621                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7651237942621 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7651237942621

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7651237942622                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7651237942622 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7651237942622

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765123794260                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765123794260 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765123794260

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765123794261                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765123794261 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765123794261

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765123794262                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765123794262 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765123794262

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765123794263                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765123794263 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765123794263

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic 17 11 13 14 16 9 10 12 15 19
+ 1 3 5 7 18
** N=39 EP=15 FDC=56
X0 1 M4_M3_CDNS_765123794260 $T=80 5580 0 0 $X=0 $Y=5190
X1 2 M4_M3_CDNS_765123794260 $T=1540 7840 0 0 $X=1460 $Y=7450
X2 3 M4_M3_CDNS_765123794260 $T=2130 6050 0 0 $X=2050 $Y=5660
X3 2 M4_M3_CDNS_765123794260 $T=2470 1570 0 0 $X=2390 $Y=1180
X4 4 M4_M3_CDNS_765123794260 $T=5260 7840 0 0 $X=5180 $Y=7450
X5 4 M4_M3_CDNS_765123794260 $T=6450 7840 0 0 $X=6370 $Y=7450
X6 4 M4_M3_CDNS_765123794260 $T=6860 1570 0 0 $X=6780 $Y=1180
X7 5 M4_M3_CDNS_765123794260 $T=7710 6520 0 0 $X=7630 $Y=6130
X8 4 M4_M3_CDNS_765123794260 $T=8050 1570 0 0 $X=7970 $Y=1180
X9 6 M4_M3_CDNS_765123794260 $T=10840 7840 0 0 $X=10760 $Y=7450
X10 6 M4_M3_CDNS_765123794260 $T=12030 7840 0 0 $X=11950 $Y=7450
X11 6 M4_M3_CDNS_765123794260 $T=12960 7840 0 0 $X=12880 $Y=7450
X12 6 M4_M3_CDNS_765123794260 $T=13370 1570 0 0 $X=13290 $Y=1180
X13 6 M4_M3_CDNS_765123794260 $T=14300 1570 0 0 $X=14220 $Y=1180
X14 6 M4_M3_CDNS_765123794260 $T=15490 1570 0 0 $X=15410 $Y=1180
X15 7 M4_M3_CDNS_765123794260 $T=16080 6990 0 0 $X=16000 $Y=6600
X16 8 M4_M3_CDNS_765123794260 $T=18280 7840 0 0 $X=18200 $Y=7450
X17 8 M4_M3_CDNS_765123794260 $T=19470 7840 0 0 $X=19390 $Y=7450
X18 8 M4_M3_CDNS_765123794260 $T=20400 7840 0 0 $X=20320 $Y=7450
X19 8 M4_M3_CDNS_765123794260 $T=21330 7840 0 0 $X=21250 $Y=7450
X20 8 M4_M3_CDNS_765123794260 $T=21740 1570 0 0 $X=21660 $Y=1180
X21 8 M4_M3_CDNS_765123794260 $T=22670 1570 0 0 $X=22590 $Y=1180
X22 8 M4_M3_CDNS_765123794260 $T=23600 1570 0 0 $X=23520 $Y=1180
X23 8 M4_M3_CDNS_765123794260 $T=24790 1570 0 0 $X=24710 $Y=1180
X24 2 M7_M6_CDNS_765123794261 $T=1540 7840 0 0 $X=1460 $Y=7450
X25 2 M7_M6_CDNS_765123794261 $T=2470 1570 0 0 $X=2390 $Y=1180
X26 4 M7_M6_CDNS_765123794261 $T=5260 7840 0 0 $X=5180 $Y=7450
X27 4 M7_M6_CDNS_765123794261 $T=6450 7840 0 0 $X=6370 $Y=7450
X28 4 M7_M6_CDNS_765123794261 $T=6860 1570 0 0 $X=6780 $Y=1180
X29 4 M7_M6_CDNS_765123794261 $T=8050 1570 0 0 $X=7970 $Y=1180
X30 6 M7_M6_CDNS_765123794261 $T=10840 7840 0 0 $X=10760 $Y=7450
X31 6 M7_M6_CDNS_765123794261 $T=12030 7840 0 0 $X=11950 $Y=7450
X32 6 M7_M6_CDNS_765123794261 $T=12960 7840 0 0 $X=12880 $Y=7450
X33 6 M7_M6_CDNS_765123794261 $T=13370 1570 0 0 $X=13290 $Y=1180
X34 6 M7_M6_CDNS_765123794261 $T=14300 1570 0 0 $X=14220 $Y=1180
X35 6 M7_M6_CDNS_765123794261 $T=15490 1570 0 0 $X=15410 $Y=1180
X36 8 M7_M6_CDNS_765123794261 $T=18280 7840 0 0 $X=18200 $Y=7450
X37 8 M7_M6_CDNS_765123794261 $T=19470 7840 0 0 $X=19390 $Y=7450
X38 8 M7_M6_CDNS_765123794261 $T=20400 7840 0 0 $X=20320 $Y=7450
X39 8 M7_M6_CDNS_765123794261 $T=21330 7840 0 0 $X=21250 $Y=7450
X40 8 M7_M6_CDNS_765123794261 $T=21740 1570 0 0 $X=21660 $Y=1180
X41 8 M7_M6_CDNS_765123794261 $T=22670 1570 0 0 $X=22590 $Y=1180
X42 8 M7_M6_CDNS_765123794261 $T=23600 1570 0 0 $X=23520 $Y=1180
X43 8 M7_M6_CDNS_765123794261 $T=24790 1570 0 0 $X=24710 $Y=1180
X44 2 M1_PO_CDNS_765123794262 $T=3580 4500 0 0 $X=3340 $Y=4250
X45 4 M1_PO_CDNS_765123794262 $T=9160 4500 0 0 $X=8920 $Y=4250
X46 6 M1_PO_CDNS_765123794262 $T=16600 4500 0 0 $X=16360 $Y=4250
X47 2 M5_M4_CDNS_765123794263 $T=3580 4500 0 0 $X=3360 $Y=4250
X48 4 M5_M4_CDNS_765123794263 $T=9160 4500 0 0 $X=8940 $Y=4250
X49 6 M5_M4_CDNS_765123794263 $T=16600 4500 0 0 $X=16380 $Y=4250
X50 8 M5_M4_CDNS_765123794263 $T=25900 4500 0 0 $X=25680 $Y=4250
X51 2 M4_M3_CDNS_765123794264 $T=3580 4500 0 0 $X=3360 $Y=4250
X52 4 M4_M3_CDNS_765123794264 $T=9160 4500 0 0 $X=8940 $Y=4250
X53 6 M4_M3_CDNS_765123794264 $T=16600 4500 0 0 $X=16380 $Y=4250
X54 8 M4_M3_CDNS_765123794264 $T=25900 4500 0 0 $X=25680 $Y=4250
X55 2 M6_M5_CDNS_765123794265 $T=3580 4500 0 0 $X=3360 $Y=4250
X56 4 M6_M5_CDNS_765123794265 $T=9160 4500 0 0 $X=8940 $Y=4250
X57 6 M6_M5_CDNS_765123794265 $T=16600 4500 0 0 $X=16380 $Y=4250
X58 8 M6_M5_CDNS_765123794265 $T=25900 4500 0 0 $X=25680 $Y=4250
X59 9 M3_M2_CDNS_765123794266 $T=610 4030 0 0 $X=530 $Y=3780
X60 1 M3_M2_CDNS_765123794266 $T=930 5440 0 0 $X=850 $Y=5190
X61 9 M3_M2_CDNS_765123794266 $T=2790 4030 0 0 $X=2710 $Y=3780
X62 10 M3_M2_CDNS_765123794266 $T=3110 3560 0 0 $X=3030 $Y=3310
X63 11 M3_M2_CDNS_765123794266 $T=4110 1490 0 0 $X=4030 $Y=1240
X64 1 M3_M2_CDNS_765123794266 $T=5580 5440 0 0 $X=5500 $Y=5190
X65 9 M3_M2_CDNS_765123794266 $T=7440 4030 0 0 $X=7360 $Y=3780
X66 12 M3_M2_CDNS_765123794266 $T=8700 3090 0 0 $X=8620 $Y=2840
X67 13 M3_M2_CDNS_765123794266 $T=9690 1490 0 0 $X=9610 $Y=1240
X68 5 M3_M2_CDNS_765123794266 $T=10230 6380 0 0 $X=10150 $Y=6130
X69 1 M3_M2_CDNS_765123794266 $T=12090 5440 0 0 $X=12010 $Y=5190
X70 9 M3_M2_CDNS_765123794266 $T=13950 4030 0 0 $X=13870 $Y=3780
X71 12 M3_M2_CDNS_765123794266 $T=15810 3090 0 0 $X=15730 $Y=2840
X72 14 M3_M2_CDNS_765123794266 $T=17130 1490 0 0 $X=17050 $Y=1240
X73 15 M3_M2_CDNS_765123794266 $T=17490 2630 0 0 $X=17410 $Y=2380
X74 5 M3_M2_CDNS_765123794266 $T=18600 6380 0 0 $X=18520 $Y=6130
X75 1 M3_M2_CDNS_765123794266 $T=20460 5440 0 0 $X=20380 $Y=5190
X76 9 M3_M2_CDNS_765123794266 $T=22320 4030 0 0 $X=22240 $Y=3780
X77 12 M3_M2_CDNS_765123794266 $T=24180 3090 0 0 $X=24100 $Y=2840
X78 16 M3_M2_CDNS_765123794266 $T=26430 1490 0 0 $X=26350 $Y=1240
X79 9 M4_M3_CDNS_765123794267 $T=610 4030 0 0 $X=530 $Y=3780
X80 1 M4_M3_CDNS_765123794267 $T=930 5440 0 0 $X=850 $Y=5190
X81 9 M4_M3_CDNS_765123794267 $T=2790 4030 0 0 $X=2710 $Y=3780
X82 1 M4_M3_CDNS_765123794267 $T=5580 5440 0 0 $X=5500 $Y=5190
X83 9 M4_M3_CDNS_765123794267 $T=7440 4030 0 0 $X=7360 $Y=3780
X84 12 M4_M3_CDNS_765123794267 $T=8700 3090 0 0 $X=8620 $Y=2840
X85 5 M4_M3_CDNS_765123794267 $T=10230 6380 0 0 $X=10150 $Y=6130
X86 1 M4_M3_CDNS_765123794267 $T=12090 5440 0 0 $X=12010 $Y=5190
X87 9 M4_M3_CDNS_765123794267 $T=13950 4030 0 0 $X=13870 $Y=3780
X88 12 M4_M3_CDNS_765123794267 $T=15810 3090 0 0 $X=15730 $Y=2840
X89 5 M4_M3_CDNS_765123794267 $T=18600 6380 0 0 $X=18520 $Y=6130
X90 1 M4_M3_CDNS_765123794267 $T=20460 5440 0 0 $X=20380 $Y=5190
X91 9 M4_M3_CDNS_765123794267 $T=22320 4030 0 0 $X=22240 $Y=3780
X92 12 M4_M3_CDNS_765123794267 $T=24180 3090 0 0 $X=24100 $Y=2840
X93 9 M5_M4_CDNS_765123794268 $T=610 4030 0 0 $X=530 $Y=3780
X94 1 M5_M4_CDNS_765123794268 $T=930 5440 0 0 $X=850 $Y=5190
X95 9 M5_M4_CDNS_765123794268 $T=2790 4030 0 0 $X=2710 $Y=3780
X96 1 M5_M4_CDNS_765123794268 $T=5580 5440 0 0 $X=5500 $Y=5190
X97 9 M5_M4_CDNS_765123794268 $T=7440 4030 0 0 $X=7360 $Y=3780
X98 12 M5_M4_CDNS_765123794268 $T=8700 3090 0 0 $X=8620 $Y=2840
X99 5 M5_M4_CDNS_765123794268 $T=10230 6380 0 0 $X=10150 $Y=6130
X100 1 M5_M4_CDNS_765123794268 $T=12090 5440 0 0 $X=12010 $Y=5190
X101 9 M5_M4_CDNS_765123794268 $T=13950 4030 0 0 $X=13870 $Y=3780
X102 12 M5_M4_CDNS_765123794268 $T=15810 3090 0 0 $X=15730 $Y=2840
X103 5 M5_M4_CDNS_765123794268 $T=18600 6380 0 0 $X=18520 $Y=6130
X104 1 M5_M4_CDNS_765123794268 $T=20460 5440 0 0 $X=20380 $Y=5190
X105 9 M5_M4_CDNS_765123794268 $T=22320 4030 0 0 $X=22240 $Y=3780
X106 12 M5_M4_CDNS_765123794268 $T=24180 3090 0 0 $X=24100 $Y=2840
X107 1 M1_PO_CDNS_765123794269 $T=930 5440 0 0 $X=830 $Y=5190
X108 17 M1_PO_CDNS_765123794269 $T=1860 4970 0 0 $X=1760 $Y=4720
X109 9 M1_PO_CDNS_765123794269 $T=2790 4030 0 0 $X=2690 $Y=3780
X110 3 M1_PO_CDNS_765123794269 $T=4650 5910 0 0 $X=4550 $Y=5660
X111 1 M1_PO_CDNS_765123794269 $T=5580 5440 0 0 $X=5480 $Y=5190
X112 17 M1_PO_CDNS_765123794269 $T=6510 4970 0 0 $X=6410 $Y=4720
X113 9 M1_PO_CDNS_765123794269 $T=7440 4030 0 0 $X=7340 $Y=3780
X114 10 M1_PO_CDNS_765123794269 $T=8370 3560 0 0 $X=8270 $Y=3310
X115 5 M1_PO_CDNS_765123794269 $T=10230 6380 0 0 $X=10130 $Y=6130
X116 3 M1_PO_CDNS_765123794269 $T=11160 5910 0 0 $X=11060 $Y=5660
X117 1 M1_PO_CDNS_765123794269 $T=12090 5440 0 0 $X=11990 $Y=5190
X118 17 M1_PO_CDNS_765123794269 $T=13020 4970 0 0 $X=12920 $Y=4720
X119 9 M1_PO_CDNS_765123794269 $T=13950 4030 0 0 $X=13850 $Y=3780
X120 10 M1_PO_CDNS_765123794269 $T=14880 3560 0 0 $X=14780 $Y=3310
X121 12 M1_PO_CDNS_765123794269 $T=15810 3090 0 0 $X=15710 $Y=2840
X122 7 M1_PO_CDNS_765123794269 $T=17670 6850 0 0 $X=17570 $Y=6600
X123 5 M1_PO_CDNS_765123794269 $T=18600 6380 0 0 $X=18500 $Y=6130
X124 3 M1_PO_CDNS_765123794269 $T=19530 5910 0 0 $X=19430 $Y=5660
X125 1 M1_PO_CDNS_765123794269 $T=20460 5440 0 0 $X=20360 $Y=5190
X126 17 M1_PO_CDNS_765123794269 $T=21390 4970 0 0 $X=21290 $Y=4720
X127 9 M1_PO_CDNS_765123794269 $T=22320 4030 0 0 $X=22220 $Y=3780
X128 10 M1_PO_CDNS_765123794269 $T=23250 3560 0 0 $X=23150 $Y=3310
X129 12 M1_PO_CDNS_765123794269 $T=24180 3090 0 0 $X=24080 $Y=2840
X130 15 M1_PO_CDNS_765123794269 $T=25110 2620 0 0 $X=25010 $Y=2370
X131 9 M2_M1_CDNS_7651237942610 $T=610 4030 0 0 $X=530 $Y=3780
X132 1 M2_M1_CDNS_7651237942610 $T=930 5440 0 0 $X=850 $Y=5190
X133 17 M2_M1_CDNS_7651237942610 $T=1860 4970 0 0 $X=1780 $Y=4720
X134 9 M2_M1_CDNS_7651237942610 $T=2790 4030 0 0 $X=2710 $Y=3780
X135 10 M2_M1_CDNS_7651237942610 $T=3110 3560 0 0 $X=3030 $Y=3310
X136 11 M2_M1_CDNS_7651237942610 $T=4110 1490 0 0 $X=4030 $Y=1240
X137 3 M2_M1_CDNS_7651237942610 $T=4650 5910 0 0 $X=4570 $Y=5660
X138 1 M2_M1_CDNS_7651237942610 $T=5580 5440 0 0 $X=5500 $Y=5190
X139 17 M2_M1_CDNS_7651237942610 $T=6510 4970 0 0 $X=6430 $Y=4720
X140 9 M2_M1_CDNS_7651237942610 $T=7440 4030 0 0 $X=7360 $Y=3780
X141 10 M2_M1_CDNS_7651237942610 $T=8370 3560 0 0 $X=8290 $Y=3310
X142 12 M2_M1_CDNS_7651237942610 $T=8700 3090 0 0 $X=8620 $Y=2840
X143 13 M2_M1_CDNS_7651237942610 $T=9690 1490 0 0 $X=9610 $Y=1240
X144 5 M2_M1_CDNS_7651237942610 $T=10230 6380 0 0 $X=10150 $Y=6130
X145 3 M2_M1_CDNS_7651237942610 $T=11160 5910 0 0 $X=11080 $Y=5660
X146 1 M2_M1_CDNS_7651237942610 $T=12090 5440 0 0 $X=12010 $Y=5190
X147 17 M2_M1_CDNS_7651237942610 $T=13020 4970 0 0 $X=12940 $Y=4720
X148 9 M2_M1_CDNS_7651237942610 $T=13950 4030 0 0 $X=13870 $Y=3780
X149 10 M2_M1_CDNS_7651237942610 $T=14880 3560 0 0 $X=14800 $Y=3310
X150 12 M2_M1_CDNS_7651237942610 $T=15810 3090 0 0 $X=15730 $Y=2840
X151 14 M2_M1_CDNS_7651237942610 $T=17130 1490 0 0 $X=17050 $Y=1240
X152 15 M2_M1_CDNS_7651237942610 $T=17490 2630 0 0 $X=17410 $Y=2380
X153 7 M2_M1_CDNS_7651237942610 $T=17670 6850 0 0 $X=17590 $Y=6600
X154 5 M2_M1_CDNS_7651237942610 $T=18600 6380 0 0 $X=18520 $Y=6130
X155 3 M2_M1_CDNS_7651237942610 $T=19530 5910 0 0 $X=19450 $Y=5660
X156 1 M2_M1_CDNS_7651237942610 $T=20460 5440 0 0 $X=20380 $Y=5190
X157 17 M2_M1_CDNS_7651237942610 $T=21390 4970 0 0 $X=21310 $Y=4720
X158 9 M2_M1_CDNS_7651237942610 $T=22320 4030 0 0 $X=22240 $Y=3780
X159 10 M2_M1_CDNS_7651237942610 $T=23250 3560 0 0 $X=23170 $Y=3310
X160 12 M2_M1_CDNS_7651237942610 $T=24180 3090 0 0 $X=24100 $Y=2840
X161 15 M2_M1_CDNS_7651237942610 $T=25110 2620 0 0 $X=25030 $Y=2370
X162 16 M2_M1_CDNS_7651237942610 $T=26430 1490 0 0 $X=26350 $Y=1240
X163 17 M3_M2_CDNS_7651237942611 $T=250 4970 0 270 $X=0 $Y=4890
X164 17 M3_M2_CDNS_7651237942611 $T=1860 4970 0 0 $X=1780 $Y=4720
X165 3 M3_M2_CDNS_7651237942611 $T=4650 5910 0 0 $X=4570 $Y=5660
X166 17 M3_M2_CDNS_7651237942611 $T=6510 4970 0 0 $X=6430 $Y=4720
X167 10 M3_M2_CDNS_7651237942611 $T=8370 3560 0 0 $X=8290 $Y=3310
X168 3 M3_M2_CDNS_7651237942611 $T=11160 5910 0 0 $X=11080 $Y=5660
X169 17 M3_M2_CDNS_7651237942611 $T=13020 4970 0 0 $X=12940 $Y=4720
X170 10 M3_M2_CDNS_7651237942611 $T=14880 3560 0 0 $X=14800 $Y=3310
X171 7 M3_M2_CDNS_7651237942611 $T=17670 6850 0 0 $X=17590 $Y=6600
X172 3 M3_M2_CDNS_7651237942611 $T=19530 5910 0 0 $X=19450 $Y=5660
X173 17 M3_M2_CDNS_7651237942611 $T=21390 4970 0 0 $X=21310 $Y=4720
X174 10 M3_M2_CDNS_7651237942611 $T=23250 3560 0 0 $X=23170 $Y=3310
X175 15 M3_M2_CDNS_7651237942611 $T=25110 2620 0 0 $X=25030 $Y=2370
X176 10 M4_M3_CDNS_7651237942614 $T=3110 3560 0 0 $X=3030 $Y=3310
X177 11 M4_M3_CDNS_7651237942614 $T=4110 1490 0 0 $X=4030 $Y=1240
X178 13 M4_M3_CDNS_7651237942614 $T=9690 1490 0 0 $X=9610 $Y=1240
X179 14 M4_M3_CDNS_7651237942614 $T=17130 1490 0 0 $X=17050 $Y=1240
X180 15 M4_M3_CDNS_7651237942614 $T=17490 2630 0 0 $X=17410 $Y=2380
X181 16 M4_M3_CDNS_7651237942614 $T=26430 1490 0 0 $X=26350 $Y=1240
X182 1 M2_M1_CDNS_7651237942615 $T=80 5580 0 0 $X=0 $Y=5190
X183 2 M2_M1_CDNS_7651237942615 $T=1540 7840 0 0 $X=1460 $Y=7450
X184 3 M2_M1_CDNS_7651237942615 $T=2130 6050 0 0 $X=2050 $Y=5660
X185 2 M2_M1_CDNS_7651237942615 $T=2470 1570 0 0 $X=2390 $Y=1180
X186 4 M2_M1_CDNS_7651237942615 $T=5260 7840 0 0 $X=5180 $Y=7450
X187 4 M2_M1_CDNS_7651237942615 $T=6450 7840 0 0 $X=6370 $Y=7450
X188 4 M2_M1_CDNS_7651237942615 $T=6860 1570 0 0 $X=6780 $Y=1180
X189 5 M2_M1_CDNS_7651237942615 $T=7710 6520 0 0 $X=7630 $Y=6130
X190 4 M2_M1_CDNS_7651237942615 $T=8050 1570 0 0 $X=7970 $Y=1180
X191 6 M2_M1_CDNS_7651237942615 $T=10840 7840 0 0 $X=10760 $Y=7450
X192 6 M2_M1_CDNS_7651237942615 $T=12030 7840 0 0 $X=11950 $Y=7450
X193 6 M2_M1_CDNS_7651237942615 $T=12960 7840 0 0 $X=12880 $Y=7450
X194 6 M2_M1_CDNS_7651237942615 $T=13370 1570 0 0 $X=13290 $Y=1180
X195 6 M2_M1_CDNS_7651237942615 $T=14300 1570 0 0 $X=14220 $Y=1180
X196 6 M2_M1_CDNS_7651237942615 $T=15490 1570 0 0 $X=15410 $Y=1180
X197 7 M2_M1_CDNS_7651237942615 $T=16080 6990 0 0 $X=16000 $Y=6600
X198 8 M2_M1_CDNS_7651237942615 $T=18280 7840 0 0 $X=18200 $Y=7450
X199 8 M2_M1_CDNS_7651237942615 $T=19470 7840 0 0 $X=19390 $Y=7450
X200 8 M2_M1_CDNS_7651237942615 $T=20400 7840 0 0 $X=20320 $Y=7450
X201 8 M2_M1_CDNS_7651237942615 $T=21330 7840 0 0 $X=21250 $Y=7450
X202 8 M2_M1_CDNS_7651237942615 $T=21740 1570 0 0 $X=21660 $Y=1180
X203 8 M2_M1_CDNS_7651237942615 $T=22670 1570 0 0 $X=22590 $Y=1180
X204 8 M2_M1_CDNS_7651237942615 $T=23600 1570 0 0 $X=23520 $Y=1180
X205 8 M2_M1_CDNS_7651237942615 $T=24790 1570 0 0 $X=24710 $Y=1180
X206 2 M2_M1_CDNS_7651237942616 $T=3580 4500 0 0 $X=3360 $Y=4250
X207 4 M2_M1_CDNS_7651237942616 $T=9160 4500 0 0 $X=8940 $Y=4250
X208 6 M2_M1_CDNS_7651237942616 $T=16600 4500 0 0 $X=16380 $Y=4250
X209 8 M2_M1_CDNS_7651237942616 $T=25900 4500 0 0 $X=25680 $Y=4250
X210 2 M3_M2_CDNS_7651237942617 $T=3580 4500 0 0 $X=3360 $Y=4250
X211 4 M3_M2_CDNS_7651237942617 $T=9160 4500 0 0 $X=8940 $Y=4250
X212 6 M3_M2_CDNS_7651237942617 $T=16600 4500 0 0 $X=16380 $Y=4250
X213 8 M3_M2_CDNS_7651237942617 $T=25900 4500 0 0 $X=25680 $Y=4250
X214 2 M7_M6_CDNS_7651237942618 $T=3580 4500 0 0 $X=3360 $Y=4250
X215 4 M7_M6_CDNS_7651237942618 $T=9160 4500 0 0 $X=8940 $Y=4250
X216 6 M7_M6_CDNS_7651237942618 $T=16600 4500 0 0 $X=16380 $Y=4250
X217 8 M7_M6_CDNS_7651237942618 $T=25900 4500 0 0 $X=25680 $Y=4250
X218 2 M6_M5_CDNS_7651237942619 $T=1540 7840 0 0 $X=1460 $Y=7450
X219 2 M6_M5_CDNS_7651237942619 $T=2470 1570 0 0 $X=2390 $Y=1180
X220 4 M6_M5_CDNS_7651237942619 $T=5260 7840 0 0 $X=5180 $Y=7450
X221 4 M6_M5_CDNS_7651237942619 $T=6450 7840 0 0 $X=6370 $Y=7450
X222 4 M6_M5_CDNS_7651237942619 $T=6860 1570 0 0 $X=6780 $Y=1180
X223 4 M6_M5_CDNS_7651237942619 $T=8050 1570 0 0 $X=7970 $Y=1180
X224 6 M6_M5_CDNS_7651237942619 $T=10840 7840 0 0 $X=10760 $Y=7450
X225 6 M6_M5_CDNS_7651237942619 $T=12030 7840 0 0 $X=11950 $Y=7450
X226 6 M6_M5_CDNS_7651237942619 $T=12960 7840 0 0 $X=12880 $Y=7450
X227 6 M6_M5_CDNS_7651237942619 $T=13370 1570 0 0 $X=13290 $Y=1180
X228 6 M6_M5_CDNS_7651237942619 $T=14300 1570 0 0 $X=14220 $Y=1180
X229 6 M6_M5_CDNS_7651237942619 $T=15490 1570 0 0 $X=15410 $Y=1180
X230 8 M6_M5_CDNS_7651237942619 $T=18280 7840 0 0 $X=18200 $Y=7450
X231 8 M6_M5_CDNS_7651237942619 $T=19470 7840 0 0 $X=19390 $Y=7450
X232 8 M6_M5_CDNS_7651237942619 $T=20400 7840 0 0 $X=20320 $Y=7450
X233 8 M6_M5_CDNS_7651237942619 $T=21330 7840 0 0 $X=21250 $Y=7450
X234 8 M6_M5_CDNS_7651237942619 $T=21740 1570 0 0 $X=21660 $Y=1180
X235 8 M6_M5_CDNS_7651237942619 $T=22670 1570 0 0 $X=22590 $Y=1180
X236 8 M6_M5_CDNS_7651237942619 $T=23600 1570 0 0 $X=23520 $Y=1180
X237 8 M6_M5_CDNS_7651237942619 $T=24790 1570 0 0 $X=24710 $Y=1180
X238 1 M6_M5_CDNS_7651237942620 $T=80 5580 0 0 $X=0 $Y=5190
X239 3 M6_M5_CDNS_7651237942620 $T=2130 6050 0 0 $X=2050 $Y=5660
X240 5 M6_M5_CDNS_7651237942620 $T=7710 6520 0 0 $X=7630 $Y=6130
X241 7 M6_M5_CDNS_7651237942620 $T=16080 6990 0 0 $X=16000 $Y=6600
X242 1 M3_M2_CDNS_7651237942621 $T=80 5580 0 0 $X=0 $Y=5190
X243 2 M3_M2_CDNS_7651237942621 $T=1540 7840 0 0 $X=1460 $Y=7450
X244 3 M3_M2_CDNS_7651237942621 $T=2130 6050 0 0 $X=2050 $Y=5660
X245 2 M3_M2_CDNS_7651237942621 $T=2470 1570 0 0 $X=2390 $Y=1180
X246 4 M3_M2_CDNS_7651237942621 $T=5260 7840 0 0 $X=5180 $Y=7450
X247 4 M3_M2_CDNS_7651237942621 $T=6450 7840 0 0 $X=6370 $Y=7450
X248 4 M3_M2_CDNS_7651237942621 $T=6860 1570 0 0 $X=6780 $Y=1180
X249 5 M3_M2_CDNS_7651237942621 $T=7710 6520 0 0 $X=7630 $Y=6130
X250 4 M3_M2_CDNS_7651237942621 $T=8050 1570 0 0 $X=7970 $Y=1180
X251 6 M3_M2_CDNS_7651237942621 $T=10840 7840 0 0 $X=10760 $Y=7450
X252 6 M3_M2_CDNS_7651237942621 $T=12030 7840 0 0 $X=11950 $Y=7450
X253 6 M3_M2_CDNS_7651237942621 $T=12960 7840 0 0 $X=12880 $Y=7450
X254 6 M3_M2_CDNS_7651237942621 $T=13370 1570 0 0 $X=13290 $Y=1180
X255 6 M3_M2_CDNS_7651237942621 $T=14300 1570 0 0 $X=14220 $Y=1180
X256 6 M3_M2_CDNS_7651237942621 $T=15490 1570 0 0 $X=15410 $Y=1180
X257 7 M3_M2_CDNS_7651237942621 $T=16080 6990 0 0 $X=16000 $Y=6600
X258 8 M3_M2_CDNS_7651237942621 $T=18280 7840 0 0 $X=18200 $Y=7450
X259 8 M3_M2_CDNS_7651237942621 $T=19470 7840 0 0 $X=19390 $Y=7450
X260 8 M3_M2_CDNS_7651237942621 $T=20400 7840 0 0 $X=20320 $Y=7450
X261 8 M3_M2_CDNS_7651237942621 $T=21330 7840 0 0 $X=21250 $Y=7450
X262 8 M3_M2_CDNS_7651237942621 $T=21740 1570 0 0 $X=21660 $Y=1180
X263 8 M3_M2_CDNS_7651237942621 $T=22670 1570 0 0 $X=22590 $Y=1180
X264 8 M3_M2_CDNS_7651237942621 $T=23600 1570 0 0 $X=23520 $Y=1180
X265 8 M3_M2_CDNS_7651237942621 $T=24790 1570 0 0 $X=24710 $Y=1180
X266 1 M5_M4_CDNS_7651237942622 $T=80 5580 0 0 $X=0 $Y=5190
X267 2 M5_M4_CDNS_7651237942622 $T=1540 7840 0 0 $X=1460 $Y=7450
X268 3 M5_M4_CDNS_7651237942622 $T=2130 6050 0 0 $X=2050 $Y=5660
X269 2 M5_M4_CDNS_7651237942622 $T=2470 1570 0 0 $X=2390 $Y=1180
X270 4 M5_M4_CDNS_7651237942622 $T=5260 7840 0 0 $X=5180 $Y=7450
X271 4 M5_M4_CDNS_7651237942622 $T=6450 7840 0 0 $X=6370 $Y=7450
X272 4 M5_M4_CDNS_7651237942622 $T=6860 1570 0 0 $X=6780 $Y=1180
X273 5 M5_M4_CDNS_7651237942622 $T=7710 6520 0 0 $X=7630 $Y=6130
X274 4 M5_M4_CDNS_7651237942622 $T=8050 1570 0 0 $X=7970 $Y=1180
X275 6 M5_M4_CDNS_7651237942622 $T=10840 7840 0 0 $X=10760 $Y=7450
X276 6 M5_M4_CDNS_7651237942622 $T=12030 7840 0 0 $X=11950 $Y=7450
X277 6 M5_M4_CDNS_7651237942622 $T=12960 7840 0 0 $X=12880 $Y=7450
X278 6 M5_M4_CDNS_7651237942622 $T=13370 1570 0 0 $X=13290 $Y=1180
X279 6 M5_M4_CDNS_7651237942622 $T=14300 1570 0 0 $X=14220 $Y=1180
X280 6 M5_M4_CDNS_7651237942622 $T=15490 1570 0 0 $X=15410 $Y=1180
X281 7 M5_M4_CDNS_7651237942622 $T=16080 6990 0 0 $X=16000 $Y=6600
X282 8 M5_M4_CDNS_7651237942622 $T=18280 7840 0 0 $X=18200 $Y=7450
X283 8 M5_M4_CDNS_7651237942622 $T=19470 7840 0 0 $X=19390 $Y=7450
X284 8 M5_M4_CDNS_7651237942622 $T=20400 7840 0 0 $X=20320 $Y=7450
X285 8 M5_M4_CDNS_7651237942622 $T=21330 7840 0 0 $X=21250 $Y=7450
X286 8 M5_M4_CDNS_7651237942622 $T=21740 1570 0 0 $X=21660 $Y=1180
X287 8 M5_M4_CDNS_7651237942622 $T=22670 1570 0 0 $X=22590 $Y=1180
X288 8 M5_M4_CDNS_7651237942622 $T=23600 1570 0 0 $X=23520 $Y=1180
X289 8 M5_M4_CDNS_7651237942622 $T=24790 1570 0 0 $X=24710 $Y=1180
X290 18 18 1 2 19 pmos1v_CDNS_765123794260 $T=1030 8610 1 0 $X=610 $Y=8170
X291 20 18 17 2 19 pmos1v_CDNS_765123794260 $T=2050 8610 0 180 $X=1540 $Y=8170
X292 21 18 1 4 19 pmos1v_CDNS_765123794260 $T=5770 8610 0 180 $X=5260 $Y=8170
X293 18 18 6 14 19 pmos1v_CDNS_765123794260 $T=16840 8610 1 0 $X=16420 $Y=8170
X294 22 18 5 8 19 pmos1v_CDNS_765123794260 $T=18790 8610 0 180 $X=18280 $Y=8170
X295 23 18 17 8 19 pmos1v_CDNS_765123794260 $T=21580 8610 0 180 $X=21070 $Y=8170
X296 22 18 12 24 19 pmos1v_CDNS_765123794260 $T=24370 8610 0 180 $X=23860 $Y=8170
X297 19 19 1 25 nmos1v_CDNS_765123794261 $T=1030 800 0 0 $X=610 $Y=240
X298 25 19 17 2 nmos1v_CDNS_765123794261 $T=1960 800 0 0 $X=1540 $Y=240
X299 19 19 3 26 nmos1v_CDNS_765123794261 $T=4750 800 0 0 $X=4330 $Y=240
X300 26 19 9 4 nmos1v_CDNS_765123794261 $T=7540 800 0 0 $X=7120 $Y=240
X301 19 19 10 4 nmos1v_CDNS_765123794261 $T=8560 800 1 180 $X=8050 $Y=240
X302 19 19 4 13 nmos1v_CDNS_765123794261 $T=9400 800 0 0 $X=8980 $Y=240
X303 27 19 1 28 nmos1v_CDNS_765123794261 $T=12190 800 0 0 $X=11770 $Y=240
X304 28 19 17 6 nmos1v_CDNS_765123794261 $T=13120 800 0 0 $X=12700 $Y=240
X305 29 19 10 6 nmos1v_CDNS_765123794261 $T=14980 800 0 0 $X=14560 $Y=240
X306 19 19 12 6 nmos1v_CDNS_765123794261 $T=16000 800 1 180 $X=15490 $Y=240
X307 19 19 6 14 nmos1v_CDNS_765123794261 $T=16840 800 0 0 $X=16420 $Y=240
X308 30 19 5 31 nmos1v_CDNS_765123794261 $T=18700 800 0 0 $X=18280 $Y=240
X309 31 19 10 8 nmos1v_CDNS_765123794261 $T=23350 800 0 0 $X=22930 $Y=240
X310 19 19 8 16 nmos1v_CDNS_765123794261 $T=26140 800 0 0 $X=25720 $Y=240
X311 19 19 9 2 nmos1v_CDNS_765123794262 $T=2980 1040 0 180 $X=2470 $Y=240
X312 19 19 2 11 nmos1v_CDNS_765123794262 $T=3820 1040 1 0 $X=3400 $Y=240
X313 26 19 1 32 nmos1v_CDNS_765123794262 $T=5680 1040 1 0 $X=5260 $Y=240
X314 32 19 17 4 nmos1v_CDNS_765123794262 $T=6610 1040 1 0 $X=6190 $Y=240
X315 19 19 5 29 nmos1v_CDNS_765123794262 $T=10330 1040 1 0 $X=9910 $Y=240
X316 29 19 3 27 nmos1v_CDNS_765123794262 $T=11260 1040 1 0 $X=10840 $Y=240
X317 27 19 9 6 nmos1v_CDNS_765123794262 $T=14050 1040 1 0 $X=13630 $Y=240
X318 19 19 7 30 nmos1v_CDNS_765123794262 $T=17770 1040 1 0 $X=17350 $Y=240
X319 31 19 3 33 nmos1v_CDNS_765123794262 $T=19630 1040 1 0 $X=19210 $Y=240
X320 33 19 1 34 nmos1v_CDNS_765123794262 $T=20560 1040 1 0 $X=20140 $Y=240
X321 34 19 17 8 nmos1v_CDNS_765123794262 $T=21490 1040 1 0 $X=21070 $Y=240
X322 33 19 9 8 nmos1v_CDNS_765123794262 $T=22420 1040 1 0 $X=22000 $Y=240
X323 30 19 12 8 nmos1v_CDNS_765123794262 $T=24280 1040 1 0 $X=23860 $Y=240
X324 19 19 15 8 nmos1v_CDNS_765123794262 $T=25300 1040 0 180 $X=24790 $Y=240
X325 18 18 9 20 19 pmos1v_CDNS_765123794263 $T=2980 8370 1 180 $X=2470 $Y=8170
X326 18 18 2 11 19 pmos1v_CDNS_765123794263 $T=3820 8370 0 0 $X=3400 $Y=8170
X327 18 18 3 4 19 pmos1v_CDNS_765123794263 $T=4750 8370 0 0 $X=4330 $Y=8170
X328 35 18 17 4 19 pmos1v_CDNS_765123794263 $T=6700 8370 1 180 $X=6190 $Y=8170
X329 21 18 9 35 19 pmos1v_CDNS_765123794263 $T=7630 8370 1 180 $X=7120 $Y=8170
X330 18 18 10 21 19 pmos1v_CDNS_765123794263 $T=8560 8370 1 180 $X=8050 $Y=8170
X331 18 18 4 13 19 pmos1v_CDNS_765123794263 $T=9400 8370 0 0 $X=8980 $Y=8170
X332 18 18 5 6 19 pmos1v_CDNS_765123794263 $T=10330 8370 0 0 $X=9910 $Y=8170
X333 36 18 3 6 19 pmos1v_CDNS_765123794263 $T=11350 8370 1 180 $X=10840 $Y=8170
X334 37 18 1 6 19 pmos1v_CDNS_765123794263 $T=12280 8370 1 180 $X=11770 $Y=8170
X335 38 18 17 6 19 pmos1v_CDNS_765123794263 $T=13210 8370 1 180 $X=12700 $Y=8170
X336 37 18 9 38 19 pmos1v_CDNS_765123794263 $T=14140 8370 1 180 $X=13630 $Y=8170
X337 36 18 10 37 19 pmos1v_CDNS_765123794263 $T=15070 8370 1 180 $X=14560 $Y=8170
X338 18 18 12 36 19 pmos1v_CDNS_765123794263 $T=16000 8370 1 180 $X=15490 $Y=8170
X339 18 18 7 8 19 pmos1v_CDNS_765123794263 $T=17770 8370 0 0 $X=17350 $Y=8170
X340 24 18 3 8 19 pmos1v_CDNS_765123794263 $T=19720 8370 1 180 $X=19210 $Y=8170
X341 39 18 1 8 19 pmos1v_CDNS_765123794263 $T=20650 8370 1 180 $X=20140 $Y=8170
X342 39 18 9 23 19 pmos1v_CDNS_765123794263 $T=22510 8370 1 180 $X=22000 $Y=8170
X343 24 18 10 39 19 pmos1v_CDNS_765123794263 $T=23440 8370 1 180 $X=22930 $Y=8170
X344 18 18 15 22 19 pmos1v_CDNS_765123794263 $T=25300 8370 1 180 $X=24790 $Y=8170
X345 18 18 8 16 19 pmos1v_CDNS_765123794263 $T=26140 8370 0 0 $X=25720 $Y=8170
M0 2 1 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1030 $Y=8370 $dt=1
M1 20 17 2 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1960 $Y=8370 $dt=1
M2 18 9 20 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=2890 $Y=8370 $dt=1
M3 11 2 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=3820 $Y=8370 $dt=1
M4 4 3 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=4750 $Y=8370 $dt=1
M5 21 1 4 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=5680 $Y=8370 $dt=1
M6 35 17 4 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=6610 $Y=8370 $dt=1
M7 21 9 35 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=7540 $Y=8370 $dt=1
M8 18 10 21 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=8470 $Y=8370 $dt=1
M9 13 4 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=9400 $Y=8370 $dt=1
M10 6 5 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=10330 $Y=8370 $dt=1
M11 36 3 6 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=11260 $Y=8370 $dt=1
M12 37 1 6 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=12190 $Y=8370 $dt=1
M13 38 17 6 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=13120 $Y=8370 $dt=1
M14 37 9 38 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=14050 $Y=8370 $dt=1
M15 36 10 37 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=14980 $Y=8370 $dt=1
M16 18 12 36 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=15910 $Y=8370 $dt=1
M17 14 6 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=16840 $Y=8370 $dt=1
M18 8 7 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=17770 $Y=8370 $dt=1
M19 22 5 8 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=18700 $Y=8370 $dt=1
M20 24 3 8 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=19630 $Y=8370 $dt=1
M21 39 1 8 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=20560 $Y=8370 $dt=1
M22 23 17 8 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21490 $Y=8370 $dt=1
M23 39 9 23 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22420 $Y=8370 $dt=1
M24 24 10 39 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23350 $Y=8370 $dt=1
M25 22 12 24 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24280 $Y=8370 $dt=1
M26 18 15 22 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25210 $Y=8370 $dt=1
M27 16 8 18 18 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26140 $Y=8370 $dt=1
.ends 4bit_CLA_logic
