* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : WallaceProjectMAC                            *
* Netlisted  : Sat Dec 13 17:03:17 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765663391800                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765663391800 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765663391800

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765663391801                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765663391801 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765663391801

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765663391802                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765663391802 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765663391802

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765663391803                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765663391803 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765663391803

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765663391804                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765663391804 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765663391804

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_765663391805                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_765663391805 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_765663391805

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_765663391806                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_765663391806 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_765663391806

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765663391807                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765663391807 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765663391807

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_765663391808                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_765663391808 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_765663391808

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765663391809                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765663391809 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765663391809

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918010                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918010 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918010

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918011                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918011 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918011

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656633918012                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656633918012 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656633918012

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918013                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918013 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918013

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918014                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918014 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918014

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918017                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918017 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918017

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656633918018                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656633918018 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656633918018

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918019                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918019 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918019

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918020                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918020 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918021                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918021 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918023                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918023 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918025                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918025 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918025

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918026                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918026 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918026

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918027                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918027 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918028                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918028 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918028

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918029                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918029 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918029

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918030                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918030 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918030

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918031                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918031 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918031

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918034                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918034 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918034

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918035                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918035 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918035

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918036                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918036 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918036

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918037                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918037 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918037

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918038                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918038 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918038

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918042                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918042 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918042

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918043                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918043 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918043

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918044                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918044 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918044

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656633918045                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656633918045 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656633918045

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656633918047                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656633918047 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656633918047

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656633918049                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656633918049 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656633918049

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918050                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918050 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918050

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656633918051                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656633918051 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656633918051

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656633918052                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656633918052 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656633918052

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656633918053                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656633918053 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656633918053

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918054                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918054 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918054

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656633918063                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656633918063 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656633918063

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918064                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918064 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918064

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765663391806                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765663391806 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765663391806

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765663391807                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765663391807 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765663391807

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918066                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918066 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918066

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656633918067                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656633918067 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656633918067

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765663391808                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765663391808 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_765663391808

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765663391809                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765663391809 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765663391809

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918010                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918010 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7656633918010

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918011                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918011 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7656633918011

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918012                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918012 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656633918012

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918013                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918013 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656633918013

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918014                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918014 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656633918014

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918015                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918015 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656633918015

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918016                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918016 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656633918016

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918017                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918017 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_7656633918017

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918018                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918018 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656633918018

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=8
X0 1 M2_M1_CDNS_7656633918020 $T=2220 -7390 0 90 $X=2090 $Y=-7470
X1 1 M2_M1_CDNS_7656633918020 $T=2220 -4680 0 90 $X=2090 $Y=-4760
X2 7 M2_M1_CDNS_7656633918020 $T=4200 -2840 0 90 $X=4070 $Y=-2920
X3 8 M2_M1_CDNS_7656633918020 $T=4570 -3920 0 90 $X=4440 $Y=-4000
X4 9 M2_M1_CDNS_7656633918025 $T=1300 -5710 0 90 $X=1170 $Y=-5840
X5 9 M2_M1_CDNS_7656633918025 $T=1300 -4270 0 90 $X=1170 $Y=-4400
X6 8 M1_PO_CDNS_7656633918063 $T=2340 -4370 0 90 $X=2090 $Y=-4470
X7 8 M1_PO_CDNS_7656633918063 $T=2930 -6480 0 90 $X=2680 $Y=-6580
X8 8 M1_PO_CDNS_7656633918063 $T=2950 -5710 0 90 $X=2700 $Y=-5810
X9 4 M1_PO_CDNS_7656633918063 $T=3490 -4140 0 90 $X=3240 $Y=-4240
X10 4 M1_PO_CDNS_7656633918063 $T=3500 -3460 0 90 $X=3250 $Y=-3560
X11 8 M2_M1_CDNS_7656633918064 $T=2340 -4370 0 90 $X=2090 $Y=-4450
X12 8 M2_M1_CDNS_7656633918064 $T=2930 -6480 0 90 $X=2680 $Y=-6560
X13 8 M2_M1_CDNS_7656633918064 $T=2950 -5710 0 90 $X=2700 $Y=-5790
X14 4 M2_M1_CDNS_7656633918064 $T=3490 -4140 0 90 $X=3240 $Y=-4220
X15 4 M2_M1_CDNS_7656633918064 $T=3500 -3460 0 90 $X=3250 $Y=-3540
X16 10 M2_M1_CDNS_7656633918064 $T=5640 -5920 0 90 $X=5390 $Y=-6000
X17 10 M2_M1_CDNS_7656633918064 $T=5640 -5080 0 90 $X=5390 $Y=-5160
X18 10 M2_M1_CDNS_7656633918064 $T=5640 -4300 0 90 $X=5390 $Y=-4380
X19 6 6 4 8 2 pmos1v_CDNS_765663391806 $T=5520 -3500 0 270 $X=5320 $Y=-4010
X20 6 6 5 7 2 pmos1v_CDNS_765663391806 $T=5520 -2570 0 270 $X=5320 $Y=-3080
X21 2 2 4 8 nmos1v_CDNS_765663391807 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X22 2 2 5 7 nmos1v_CDNS_765663391807 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X23 4 M2_M1_CDNS_7656633918066 $T=3500 -4810 0 0 $X=3250 $Y=-4940
X24 4 M2_M1_CDNS_7656633918066 $T=3500 -1930 0 0 $X=3250 $Y=-2060
X25 7 M2_M1_CDNS_7656633918066 $T=4210 -6730 0 0 $X=3960 $Y=-6860
X26 7 M2_M1_CDNS_7656633918066 $T=4210 -5370 0 0 $X=3960 $Y=-5500
X27 8 M2_M1_CDNS_7656633918066 $T=4540 -5740 0 0 $X=4290 $Y=-5870
X28 5 M2_M1_CDNS_7656633918066 $T=4960 -4960 0 0 $X=4710 $Y=-5090
X29 5 M2_M1_CDNS_7656633918066 $T=4960 -2500 0 0 $X=4710 $Y=-2630
X30 4 M1_PO_CDNS_7656633918067 $T=3500 -4810 0 0 $X=3260 $Y=-4910
X31 7 M1_PO_CDNS_7656633918067 $T=4210 -6730 0 0 $X=3970 $Y=-6830
X32 7 M1_PO_CDNS_7656633918067 $T=4210 -5370 0 0 $X=3970 $Y=-5470
X33 8 M1_PO_CDNS_7656633918067 $T=4540 -5740 0 0 $X=4300 $Y=-5840
X34 5 M1_PO_CDNS_7656633918067 $T=4960 -4960 0 0 $X=4720 $Y=-5060
X35 5 M1_PO_CDNS_7656633918067 $T=4960 -2500 0 0 $X=4720 $Y=-2600
X36 1 5 10 2 6 pmos1v_CDNS_765663391808 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 2 7 3 nmos1v_CDNS_765663391809 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 10 6 7 2 pmos1v_CDNS_7656633918010 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 6 8 11 2 pmos1v_CDNS_7656633918011 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 3 7 11 2 6 pmos1v_CDNS_7656633918012 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X41 2 3 8 2 nmos1v_CDNS_7656633918013 $T=1570 -6390 0 270 $X=1370 $Y=-6840
X42 9 1 8 2 nmos1v_CDNS_7656633918013 $T=1570 -4430 0 270 $X=1370 $Y=-4880
X43 9 7 2 2 nmos1v_CDNS_7656633918014 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 4 1 12 2 nmos1v_CDNS_7656633918015 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 2 5 12 nmos1v_CDNS_7656633918016 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 10 8 6 2 pmos1v_CDNS_7656633918017 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 10 4 1 2 6 pmos1v_CDNS_7656633918018 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 2 8 3 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 2 7 9 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=6.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-5550 $dt=0
M2 9 8 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M3 2 4 8 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-3590 $dt=0
M4 2 5 7 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1580 $Y=-2660 $dt=0
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656633918057                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656633918057 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656633918057

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918058                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918058 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918058

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918059                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918059 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918059

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918060                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918060 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918060

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656633918061                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656633918061 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656633918061

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656633918062                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656633918062 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656633918062

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765663391800                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765663391800 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_765663391800

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765663391801                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765663391801 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765663391801

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765663391802                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765663391802 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_765663391802

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765663391803                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765663391803 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765663391803

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765663391804                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765663391804 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765663391804

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765663391805                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765663391805 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765663391805

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=0
X0 1 M2_M1_CDNS_7656633918020 $T=1510 -2070 0 0 $X=1430 $Y=-2200
X1 1 M2_M1_CDNS_7656633918020 $T=3010 -2070 0 0 $X=2930 $Y=-2200
X2 5 M3_M2_CDNS_7656633918027 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X3 5 M2_M1_CDNS_7656633918028 $T=5170 -2000 0 0 $X=5090 $Y=-2250
X4 2 M1_PO_CDNS_7656633918062 $T=1870 -1670 0 0 $X=1770 $Y=-1790
X5 1 M1_PO_CDNS_7656633918062 $T=2510 -2070 0 0 $X=2410 $Y=-2190
X6 6 M1_PO_CDNS_7656633918062 $T=4500 -2020 0 0 $X=4400 $Y=-2140
X7 4 5 6 nmos1v_CDNS_765663391800 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X8 3 5 6 4 pmos1v_CDNS_765663391801 $T=4560 -1510 0 0 $X=3880 $Y=-1710
X9 4 1 7 nmos1v_CDNS_765663391802 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X10 3 2 6 4 pmos1v_CDNS_765663391803 $T=1930 -1320 0 0 $X=1250 $Y=-1520
X11 3 6 1 4 pmos1v_CDNS_765663391804 $T=2430 -1320 1 180 $X=1980 $Y=-1520
X12 6 2 7 4 nmos1v_CDNS_765663391805 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR 1 2 3 4 5 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X0 6 M2_M1_CDNS_7656633918020 $T=690 3330 0 0 $X=610 $Y=3200
X1 1 M2_M1_CDNS_7656633918020 $T=1190 1490 0 0 $X=1110 $Y=1360
X2 1 M2_M1_CDNS_7656633918020 $T=2520 1490 0 0 $X=2440 $Y=1360
X3 6 M2_M1_CDNS_7656633918020 $T=2550 3330 0 0 $X=2470 $Y=3200
X4 4 M5_M4_CDNS_7656633918057 $T=1850 2810 0 90 $X=1600 $Y=2590
X5 4 M4_M3_CDNS_7656633918058 $T=1850 2810 0 90 $X=1600 $Y=2590
X6 4 M3_M2_CDNS_7656633918059 $T=1850 2810 0 90 $X=1600 $Y=2590
X7 4 M2_M1_CDNS_7656633918060 $T=1850 2810 0 90 $X=1600 $Y=2590
X8 4 M6_M5_CDNS_7656633918061 $T=1850 2810 0 90 $X=1600 $Y=2590
X9 7 M1_PO_CDNS_7656633918062 $T=2470 2570 0 0 $X=2370 $Y=2450
X10 1 M1_PO_CDNS_7656633918063 $T=320 1490 0 0 $X=220 $Y=1240
X11 5 M1_PO_CDNS_7656633918063 $T=1540 2050 0 0 $X=1440 $Y=1800
X12 5 M1_PO_CDNS_7656633918063 $T=3400 2050 0 0 $X=3300 $Y=1800
X13 1 M2_M1_CDNS_7656633918064 $T=320 1490 0 0 $X=240 $Y=1240
X14 5 M2_M1_CDNS_7656633918064 $T=1540 2050 0 0 $X=1460 $Y=1800
X15 5 M2_M1_CDNS_7656633918064 $T=3400 2050 0 0 $X=3320 $Y=1800
X16 2 2 1 6 3 pmos1v_CDNS_765663391806 $T=420 3660 0 0 $X=0 $Y=3460
X17 1 2 5 4 3 pmos1v_CDNS_765663391806 $T=1350 3660 0 0 $X=930 $Y=3460
X18 6 2 7 4 3 pmos1v_CDNS_765663391806 $T=2370 3660 1 180 $X=1860 $Y=3460
X19 2 2 5 7 3 pmos1v_CDNS_765663391806 $T=3300 3660 1 180 $X=2790 $Y=3460
X20 3 3 1 6 nmos1v_CDNS_765663391807 $T=420 800 0 0 $X=0 $Y=240
X21 4 3 5 6 nmos1v_CDNS_765663391807 $T=1440 800 1 180 $X=930 $Y=240
X22 4 3 7 1 nmos1v_CDNS_765663391807 $T=2280 800 0 0 $X=1860 $Y=240
X23 3 3 5 7 nmos1v_CDNS_765663391807 $T=3300 800 1 180 $X=2790 $Y=240
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=420 $Y=800 $dt=0
M1 4 5 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1350 $Y=800 $dt=0
M2 1 7 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=2280 $Y=800 $dt=0
M3 3 5 7 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=3210 $Y=800 $dt=0
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7656633918068                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7656633918068 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7656633918068

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656633918069                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656633918069 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656633918069

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656633918070                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656633918070 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656633918070

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656633918071                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656633918071 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656633918071

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7656633918072                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7656633918072 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7656633918072

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918074                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918074 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918074

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M7_M6_CDNS_7656633918075                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M7_M6_CDNS_7656633918075 1
** N=1 EP=1 FDC=0
.ends M7_M6_CDNS_7656633918075

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656633918076                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656633918076 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656633918076

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M6_M5_CDNS_7656633918077                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M6_M5_CDNS_7656633918077 1
** N=1 EP=1 FDC=0
.ends M6_M5_CDNS_7656633918077

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7656633918078                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7656633918078 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7656633918078

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7656633918079                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7656633918079 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7656633918079

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918019                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918019 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656633918019

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918020                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918020 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656633918020

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39
*.DEVICECLIMB
** N=39 EP=39 FDC=54
X0 2 M5_M4_CDNS_765663391808 $T=610 4030 0 0 $X=530 $Y=3780
X1 1 M5_M4_CDNS_765663391808 $T=930 5440 0 0 $X=850 $Y=5190
X2 2 M5_M4_CDNS_765663391808 $T=2790 4030 0 0 $X=2710 $Y=3780
X3 1 M5_M4_CDNS_765663391808 $T=5580 5440 0 0 $X=5500 $Y=5190
X4 2 M5_M4_CDNS_765663391808 $T=7440 4030 0 0 $X=7360 $Y=3780
X5 10 M5_M4_CDNS_765663391808 $T=8700 3090 0 0 $X=8620 $Y=2840
X6 9 M5_M4_CDNS_765663391808 $T=10230 6380 0 0 $X=10150 $Y=6130
X7 1 M5_M4_CDNS_765663391808 $T=12090 5440 0 0 $X=12010 $Y=5190
X8 2 M5_M4_CDNS_765663391808 $T=13950 4030 0 0 $X=13870 $Y=3780
X9 10 M5_M4_CDNS_765663391808 $T=15810 3090 0 0 $X=15730 $Y=2840
X10 9 M5_M4_CDNS_765663391808 $T=18600 6380 0 0 $X=18520 $Y=6130
X11 1 M5_M4_CDNS_765663391808 $T=20460 5440 0 0 $X=20380 $Y=5190
X12 2 M5_M4_CDNS_765663391808 $T=22320 4030 0 0 $X=22240 $Y=3780
X13 10 M5_M4_CDNS_765663391808 $T=24180 3090 0 0 $X=24100 $Y=2840
X14 2 M2_M1_CDNS_765663391809 $T=610 4030 0 0 $X=530 $Y=3780
X15 1 M2_M1_CDNS_765663391809 $T=930 5440 0 0 $X=850 $Y=5190
X16 3 M2_M1_CDNS_765663391809 $T=1860 4970 0 0 $X=1780 $Y=4720
X17 2 M2_M1_CDNS_765663391809 $T=2790 4030 0 0 $X=2710 $Y=3780
X18 7 M2_M1_CDNS_765663391809 $T=3110 3560 0 0 $X=3030 $Y=3310
X19 8 M2_M1_CDNS_765663391809 $T=4110 1490 0 0 $X=4030 $Y=1240
X20 6 M2_M1_CDNS_765663391809 $T=4650 5910 0 0 $X=4570 $Y=5660
X21 1 M2_M1_CDNS_765663391809 $T=5580 5440 0 0 $X=5500 $Y=5190
X22 3 M2_M1_CDNS_765663391809 $T=6510 4970 0 0 $X=6430 $Y=4720
X23 2 M2_M1_CDNS_765663391809 $T=7440 4030 0 0 $X=7360 $Y=3780
X24 7 M2_M1_CDNS_765663391809 $T=8370 3560 0 0 $X=8290 $Y=3310
X25 10 M2_M1_CDNS_765663391809 $T=8700 3090 0 0 $X=8620 $Y=2840
X26 11 M2_M1_CDNS_765663391809 $T=9690 1490 0 0 $X=9610 $Y=1240
X27 9 M2_M1_CDNS_765663391809 $T=10230 6380 0 0 $X=10150 $Y=6130
X28 6 M2_M1_CDNS_765663391809 $T=11160 5910 0 0 $X=11080 $Y=5660
X29 1 M2_M1_CDNS_765663391809 $T=12090 5440 0 0 $X=12010 $Y=5190
X30 3 M2_M1_CDNS_765663391809 $T=13020 4970 0 0 $X=12940 $Y=4720
X31 2 M2_M1_CDNS_765663391809 $T=13950 4030 0 0 $X=13870 $Y=3780
X32 7 M2_M1_CDNS_765663391809 $T=14880 3560 0 0 $X=14800 $Y=3310
X33 10 M2_M1_CDNS_765663391809 $T=15810 3090 0 0 $X=15730 $Y=2840
X34 13 M2_M1_CDNS_765663391809 $T=17130 1490 0 0 $X=17050 $Y=1240
X35 14 M2_M1_CDNS_765663391809 $T=17490 2630 0 0 $X=17410 $Y=2380
X36 12 M2_M1_CDNS_765663391809 $T=17670 6850 0 0 $X=17590 $Y=6600
X37 9 M2_M1_CDNS_765663391809 $T=18600 6380 0 0 $X=18520 $Y=6130
X38 6 M2_M1_CDNS_765663391809 $T=19530 5910 0 0 $X=19450 $Y=5660
X39 1 M2_M1_CDNS_765663391809 $T=20460 5440 0 0 $X=20380 $Y=5190
X40 3 M2_M1_CDNS_765663391809 $T=21390 4970 0 0 $X=21310 $Y=4720
X41 2 M2_M1_CDNS_765663391809 $T=22320 4030 0 0 $X=22240 $Y=3780
X42 7 M2_M1_CDNS_765663391809 $T=23250 3560 0 0 $X=23170 $Y=3310
X43 10 M2_M1_CDNS_765663391809 $T=24180 3090 0 0 $X=24100 $Y=2840
X44 14 M2_M1_CDNS_765663391809 $T=25110 2620 0 0 $X=25030 $Y=2370
X45 15 M2_M1_CDNS_765663391809 $T=26430 1490 0 0 $X=26350 $Y=1240
X46 2 M4_M3_CDNS_7656633918010 $T=610 4030 0 0 $X=530 $Y=3780
X47 1 M4_M3_CDNS_7656633918010 $T=930 5440 0 0 $X=850 $Y=5190
X48 2 M4_M3_CDNS_7656633918010 $T=2790 4030 0 0 $X=2710 $Y=3780
X49 1 M4_M3_CDNS_7656633918010 $T=5580 5440 0 0 $X=5500 $Y=5190
X50 2 M4_M3_CDNS_7656633918010 $T=7440 4030 0 0 $X=7360 $Y=3780
X51 10 M4_M3_CDNS_7656633918010 $T=8700 3090 0 0 $X=8620 $Y=2840
X52 9 M4_M3_CDNS_7656633918010 $T=10230 6380 0 0 $X=10150 $Y=6130
X53 1 M4_M3_CDNS_7656633918010 $T=12090 5440 0 0 $X=12010 $Y=5190
X54 2 M4_M3_CDNS_7656633918010 $T=13950 4030 0 0 $X=13870 $Y=3780
X55 10 M4_M3_CDNS_7656633918010 $T=15810 3090 0 0 $X=15730 $Y=2840
X56 9 M4_M3_CDNS_7656633918010 $T=18600 6380 0 0 $X=18520 $Y=6130
X57 1 M4_M3_CDNS_7656633918010 $T=20460 5440 0 0 $X=20380 $Y=5190
X58 2 M4_M3_CDNS_7656633918010 $T=22320 4030 0 0 $X=22240 $Y=3780
X59 10 M4_M3_CDNS_7656633918010 $T=24180 3090 0 0 $X=24100 $Y=2840
X60 2 M3_M2_CDNS_7656633918011 $T=610 4030 0 0 $X=530 $Y=3780
X61 1 M3_M2_CDNS_7656633918011 $T=930 5440 0 0 $X=850 $Y=5190
X62 2 M3_M2_CDNS_7656633918011 $T=2790 4030 0 0 $X=2710 $Y=3780
X63 7 M3_M2_CDNS_7656633918011 $T=3110 3560 0 0 $X=3030 $Y=3310
X64 8 M3_M2_CDNS_7656633918011 $T=4110 1490 0 0 $X=4030 $Y=1240
X65 1 M3_M2_CDNS_7656633918011 $T=5580 5440 0 0 $X=5500 $Y=5190
X66 2 M3_M2_CDNS_7656633918011 $T=7440 4030 0 0 $X=7360 $Y=3780
X67 10 M3_M2_CDNS_7656633918011 $T=8700 3090 0 0 $X=8620 $Y=2840
X68 11 M3_M2_CDNS_7656633918011 $T=9690 1490 0 0 $X=9610 $Y=1240
X69 9 M3_M2_CDNS_7656633918011 $T=10230 6380 0 0 $X=10150 $Y=6130
X70 1 M3_M2_CDNS_7656633918011 $T=12090 5440 0 0 $X=12010 $Y=5190
X71 2 M3_M2_CDNS_7656633918011 $T=13950 4030 0 0 $X=13870 $Y=3780
X72 10 M3_M2_CDNS_7656633918011 $T=15810 3090 0 0 $X=15730 $Y=2840
X73 13 M3_M2_CDNS_7656633918011 $T=17130 1490 0 0 $X=17050 $Y=1240
X74 14 M3_M2_CDNS_7656633918011 $T=17490 2630 0 0 $X=17410 $Y=2380
X75 9 M3_M2_CDNS_7656633918011 $T=18600 6380 0 0 $X=18520 $Y=6130
X76 1 M3_M2_CDNS_7656633918011 $T=20460 5440 0 0 $X=20380 $Y=5190
X77 2 M3_M2_CDNS_7656633918011 $T=22320 4030 0 0 $X=22240 $Y=3780
X78 10 M3_M2_CDNS_7656633918011 $T=24180 3090 0 0 $X=24100 $Y=2840
X79 15 M3_M2_CDNS_7656633918011 $T=26430 1490 0 0 $X=26350 $Y=1240
X80 3 M3_M2_CDNS_7656633918027 $T=250 4970 0 90 $X=0 $Y=4890
X81 3 M3_M2_CDNS_7656633918027 $T=1860 4970 0 0 $X=1780 $Y=4720
X82 6 M3_M2_CDNS_7656633918027 $T=4650 5910 0 0 $X=4570 $Y=5660
X83 3 M3_M2_CDNS_7656633918027 $T=6510 4970 0 0 $X=6430 $Y=4720
X84 7 M3_M2_CDNS_7656633918027 $T=8370 3560 0 0 $X=8290 $Y=3310
X85 6 M3_M2_CDNS_7656633918027 $T=11160 5910 0 0 $X=11080 $Y=5660
X86 3 M3_M2_CDNS_7656633918027 $T=13020 4970 0 0 $X=12940 $Y=4720
X87 7 M3_M2_CDNS_7656633918027 $T=14880 3560 0 0 $X=14800 $Y=3310
X88 12 M3_M2_CDNS_7656633918027 $T=17670 6850 0 0 $X=17590 $Y=6600
X89 6 M3_M2_CDNS_7656633918027 $T=19530 5910 0 0 $X=19450 $Y=5660
X90 3 M3_M2_CDNS_7656633918027 $T=21390 4970 0 0 $X=21310 $Y=4720
X91 7 M3_M2_CDNS_7656633918027 $T=23250 3560 0 0 $X=23170 $Y=3310
X92 14 M3_M2_CDNS_7656633918027 $T=25110 2620 0 0 $X=25030 $Y=2370
X93 3 M2_M1_CDNS_7656633918028 $T=250 4970 0 90 $X=0 $Y=4890
X94 7 M4_M3_CDNS_7656633918036 $T=3110 3560 0 0 $X=3030 $Y=3310
X95 8 M4_M3_CDNS_7656633918036 $T=4110 1490 0 0 $X=4030 $Y=1240
X96 11 M4_M3_CDNS_7656633918036 $T=9690 1490 0 0 $X=9610 $Y=1240
X97 13 M4_M3_CDNS_7656633918036 $T=17130 1490 0 0 $X=17050 $Y=1240
X98 14 M4_M3_CDNS_7656633918036 $T=17490 2630 0 0 $X=17410 $Y=2380
X99 15 M4_M3_CDNS_7656633918036 $T=26430 1490 0 0 $X=26350 $Y=1240
X100 16 M5_M4_CDNS_7656633918057 $T=3580 4500 0 0 $X=3360 $Y=4250
X101 17 M5_M4_CDNS_7656633918057 $T=9160 4500 0 0 $X=8940 $Y=4250
X102 18 M5_M4_CDNS_7656633918057 $T=16600 4500 0 0 $X=16380 $Y=4250
X103 19 M5_M4_CDNS_7656633918057 $T=25900 4500 0 0 $X=25680 $Y=4250
X104 16 M4_M3_CDNS_7656633918058 $T=3580 4500 0 0 $X=3360 $Y=4250
X105 17 M4_M3_CDNS_7656633918058 $T=9160 4500 0 0 $X=8940 $Y=4250
X106 18 M4_M3_CDNS_7656633918058 $T=16600 4500 0 0 $X=16380 $Y=4250
X107 19 M4_M3_CDNS_7656633918058 $T=25900 4500 0 0 $X=25680 $Y=4250
X108 16 M3_M2_CDNS_7656633918059 $T=3580 4500 0 0 $X=3360 $Y=4250
X109 17 M3_M2_CDNS_7656633918059 $T=9160 4500 0 0 $X=8940 $Y=4250
X110 18 M3_M2_CDNS_7656633918059 $T=16600 4500 0 0 $X=16380 $Y=4250
X111 19 M3_M2_CDNS_7656633918059 $T=25900 4500 0 0 $X=25680 $Y=4250
X112 16 M2_M1_CDNS_7656633918060 $T=3580 4500 0 0 $X=3360 $Y=4250
X113 17 M2_M1_CDNS_7656633918060 $T=9160 4500 0 0 $X=8940 $Y=4250
X114 18 M2_M1_CDNS_7656633918060 $T=16600 4500 0 0 $X=16380 $Y=4250
X115 19 M2_M1_CDNS_7656633918060 $T=25900 4500 0 0 $X=25680 $Y=4250
X116 4 4 2 20 5 pmos1v_CDNS_765663391806 $T=2980 8370 1 180 $X=2470 $Y=8170
X117 4 4 16 8 5 pmos1v_CDNS_765663391806 $T=3820 8370 0 0 $X=3400 $Y=8170
X118 4 4 6 17 5 pmos1v_CDNS_765663391806 $T=4750 8370 0 0 $X=4330 $Y=8170
X119 21 4 3 17 5 pmos1v_CDNS_765663391806 $T=6700 8370 1 180 $X=6190 $Y=8170
X120 22 4 2 21 5 pmos1v_CDNS_765663391806 $T=7630 8370 1 180 $X=7120 $Y=8170
X121 4 4 7 22 5 pmos1v_CDNS_765663391806 $T=8560 8370 1 180 $X=8050 $Y=8170
X122 4 4 17 11 5 pmos1v_CDNS_765663391806 $T=9400 8370 0 0 $X=8980 $Y=8170
X123 4 4 9 18 5 pmos1v_CDNS_765663391806 $T=10330 8370 0 0 $X=9910 $Y=8170
X124 23 4 6 18 5 pmos1v_CDNS_765663391806 $T=11350 8370 1 180 $X=10840 $Y=8170
X125 24 4 1 18 5 pmos1v_CDNS_765663391806 $T=12280 8370 1 180 $X=11770 $Y=8170
X126 25 4 3 18 5 pmos1v_CDNS_765663391806 $T=13210 8370 1 180 $X=12700 $Y=8170
X127 24 4 2 25 5 pmos1v_CDNS_765663391806 $T=14140 8370 1 180 $X=13630 $Y=8170
X128 23 4 7 24 5 pmos1v_CDNS_765663391806 $T=15070 8370 1 180 $X=14560 $Y=8170
X129 4 4 10 23 5 pmos1v_CDNS_765663391806 $T=16000 8370 1 180 $X=15490 $Y=8170
X130 4 4 12 19 5 pmos1v_CDNS_765663391806 $T=17770 8370 0 0 $X=17350 $Y=8170
X131 26 4 6 19 5 pmos1v_CDNS_765663391806 $T=19720 8370 1 180 $X=19210 $Y=8170
X132 27 4 1 19 5 pmos1v_CDNS_765663391806 $T=20650 8370 1 180 $X=20140 $Y=8170
X133 27 4 2 28 5 pmos1v_CDNS_765663391806 $T=22510 8370 1 180 $X=22000 $Y=8170
X134 26 4 7 27 5 pmos1v_CDNS_765663391806 $T=23440 8370 1 180 $X=22930 $Y=8170
X135 4 4 14 29 5 pmos1v_CDNS_765663391806 $T=25300 8370 1 180 $X=24790 $Y=8170
X136 4 4 19 15 5 pmos1v_CDNS_765663391806 $T=26140 8370 0 0 $X=25720 $Y=8170
X137 5 5 1 30 nmos1v_CDNS_765663391807 $T=1030 800 0 0 $X=610 $Y=240
X138 30 5 3 16 nmos1v_CDNS_765663391807 $T=1960 800 0 0 $X=1540 $Y=240
X139 5 5 6 31 nmos1v_CDNS_765663391807 $T=4750 800 0 0 $X=4330 $Y=240
X140 31 5 2 17 nmos1v_CDNS_765663391807 $T=7540 800 0 0 $X=7120 $Y=240
X141 5 5 7 17 nmos1v_CDNS_765663391807 $T=8560 800 1 180 $X=8050 $Y=240
X142 5 5 17 11 nmos1v_CDNS_765663391807 $T=9400 800 0 0 $X=8980 $Y=240
X143 32 5 1 33 nmos1v_CDNS_765663391807 $T=12190 800 0 0 $X=11770 $Y=240
X144 33 5 3 18 nmos1v_CDNS_765663391807 $T=13120 800 0 0 $X=12700 $Y=240
X145 34 5 7 18 nmos1v_CDNS_765663391807 $T=14980 800 0 0 $X=14560 $Y=240
X146 5 5 10 18 nmos1v_CDNS_765663391807 $T=16000 800 1 180 $X=15490 $Y=240
X147 5 5 18 13 nmos1v_CDNS_765663391807 $T=16840 800 0 0 $X=16420 $Y=240
X148 35 5 9 36 nmos1v_CDNS_765663391807 $T=18700 800 0 0 $X=18280 $Y=240
X149 36 5 7 19 nmos1v_CDNS_765663391807 $T=23350 800 0 0 $X=22930 $Y=240
X150 5 5 19 15 nmos1v_CDNS_765663391807 $T=26140 800 0 0 $X=25720 $Y=240
X151 1 M4_M3_CDNS_7656633918068 $T=80 5580 0 0 $X=0 $Y=5190
X152 16 M4_M3_CDNS_7656633918068 $T=1540 7840 0 0 $X=1460 $Y=7450
X153 6 M4_M3_CDNS_7656633918068 $T=2130 6050 0 0 $X=2050 $Y=5660
X154 16 M4_M3_CDNS_7656633918068 $T=2470 1570 0 0 $X=2390 $Y=1180
X155 17 M4_M3_CDNS_7656633918068 $T=5260 7840 0 0 $X=5180 $Y=7450
X156 17 M4_M3_CDNS_7656633918068 $T=6450 7840 0 0 $X=6370 $Y=7450
X157 17 M4_M3_CDNS_7656633918068 $T=6860 1570 0 0 $X=6780 $Y=1180
X158 9 M4_M3_CDNS_7656633918068 $T=7710 6520 0 0 $X=7630 $Y=6130
X159 17 M4_M3_CDNS_7656633918068 $T=8050 1570 0 0 $X=7970 $Y=1180
X160 18 M4_M3_CDNS_7656633918068 $T=10840 7840 0 0 $X=10760 $Y=7450
X161 18 M4_M3_CDNS_7656633918068 $T=12030 7840 0 0 $X=11950 $Y=7450
X162 18 M4_M3_CDNS_7656633918068 $T=12960 7840 0 0 $X=12880 $Y=7450
X163 18 M4_M3_CDNS_7656633918068 $T=13370 1570 0 0 $X=13290 $Y=1180
X164 18 M4_M3_CDNS_7656633918068 $T=14300 1570 0 0 $X=14220 $Y=1180
X165 18 M4_M3_CDNS_7656633918068 $T=15490 1570 0 0 $X=15410 $Y=1180
X166 12 M4_M3_CDNS_7656633918068 $T=16080 6990 0 0 $X=16000 $Y=6600
X167 19 M4_M3_CDNS_7656633918068 $T=18280 7840 0 0 $X=18200 $Y=7450
X168 19 M4_M3_CDNS_7656633918068 $T=19470 7840 0 0 $X=19390 $Y=7450
X169 19 M4_M3_CDNS_7656633918068 $T=20400 7840 0 0 $X=20320 $Y=7450
X170 19 M4_M3_CDNS_7656633918068 $T=21330 7840 0 0 $X=21250 $Y=7450
X171 19 M4_M3_CDNS_7656633918068 $T=21740 1570 0 0 $X=21660 $Y=1180
X172 19 M4_M3_CDNS_7656633918068 $T=22670 1570 0 0 $X=22590 $Y=1180
X173 19 M4_M3_CDNS_7656633918068 $T=23600 1570 0 0 $X=23520 $Y=1180
X174 19 M4_M3_CDNS_7656633918068 $T=24790 1570 0 0 $X=24710 $Y=1180
X175 16 M7_M6_CDNS_7656633918069 $T=1540 7840 0 0 $X=1460 $Y=7450
X176 16 M7_M6_CDNS_7656633918069 $T=2470 1570 0 0 $X=2390 $Y=1180
X177 17 M7_M6_CDNS_7656633918069 $T=5260 7840 0 0 $X=5180 $Y=7450
X178 17 M7_M6_CDNS_7656633918069 $T=6450 7840 0 0 $X=6370 $Y=7450
X179 17 M7_M6_CDNS_7656633918069 $T=6860 1570 0 0 $X=6780 $Y=1180
X180 17 M7_M6_CDNS_7656633918069 $T=8050 1570 0 0 $X=7970 $Y=1180
X181 18 M7_M6_CDNS_7656633918069 $T=10840 7840 0 0 $X=10760 $Y=7450
X182 18 M7_M6_CDNS_7656633918069 $T=12030 7840 0 0 $X=11950 $Y=7450
X183 18 M7_M6_CDNS_7656633918069 $T=12960 7840 0 0 $X=12880 $Y=7450
X184 18 M7_M6_CDNS_7656633918069 $T=13370 1570 0 0 $X=13290 $Y=1180
X185 18 M7_M6_CDNS_7656633918069 $T=14300 1570 0 0 $X=14220 $Y=1180
X186 18 M7_M6_CDNS_7656633918069 $T=15490 1570 0 0 $X=15410 $Y=1180
X187 19 M7_M6_CDNS_7656633918069 $T=18280 7840 0 0 $X=18200 $Y=7450
X188 19 M7_M6_CDNS_7656633918069 $T=19470 7840 0 0 $X=19390 $Y=7450
X189 19 M7_M6_CDNS_7656633918069 $T=20400 7840 0 0 $X=20320 $Y=7450
X190 19 M7_M6_CDNS_7656633918069 $T=21330 7840 0 0 $X=21250 $Y=7450
X191 19 M7_M6_CDNS_7656633918069 $T=21740 1570 0 0 $X=21660 $Y=1180
X192 19 M7_M6_CDNS_7656633918069 $T=22670 1570 0 0 $X=22590 $Y=1180
X193 19 M7_M6_CDNS_7656633918069 $T=23600 1570 0 0 $X=23520 $Y=1180
X194 19 M7_M6_CDNS_7656633918069 $T=24790 1570 0 0 $X=24710 $Y=1180
X195 16 M1_PO_CDNS_7656633918070 $T=3580 4500 0 0 $X=3340 $Y=4250
X196 17 M1_PO_CDNS_7656633918070 $T=9160 4500 0 0 $X=8920 $Y=4250
X197 18 M1_PO_CDNS_7656633918070 $T=16600 4500 0 0 $X=16360 $Y=4250
X198 16 M6_M5_CDNS_7656633918071 $T=3580 4500 0 0 $X=3360 $Y=4250
X199 17 M6_M5_CDNS_7656633918071 $T=9160 4500 0 0 $X=8940 $Y=4250
X200 18 M6_M5_CDNS_7656633918071 $T=16600 4500 0 0 $X=16380 $Y=4250
X201 19 M6_M5_CDNS_7656633918071 $T=25900 4500 0 0 $X=25680 $Y=4250
X202 1 M1_PO_CDNS_7656633918072 $T=930 5440 0 0 $X=830 $Y=5190
X203 3 M1_PO_CDNS_7656633918072 $T=1860 4970 0 0 $X=1760 $Y=4720
X204 2 M1_PO_CDNS_7656633918072 $T=2790 4030 0 0 $X=2690 $Y=3780
X205 6 M1_PO_CDNS_7656633918072 $T=4650 5910 0 0 $X=4550 $Y=5660
X206 1 M1_PO_CDNS_7656633918072 $T=5580 5440 0 0 $X=5480 $Y=5190
X207 3 M1_PO_CDNS_7656633918072 $T=6510 4970 0 0 $X=6410 $Y=4720
X208 2 M1_PO_CDNS_7656633918072 $T=7440 4030 0 0 $X=7340 $Y=3780
X209 7 M1_PO_CDNS_7656633918072 $T=8370 3560 0 0 $X=8270 $Y=3310
X210 9 M1_PO_CDNS_7656633918072 $T=10230 6380 0 0 $X=10130 $Y=6130
X211 6 M1_PO_CDNS_7656633918072 $T=11160 5910 0 0 $X=11060 $Y=5660
X212 1 M1_PO_CDNS_7656633918072 $T=12090 5440 0 0 $X=11990 $Y=5190
X213 3 M1_PO_CDNS_7656633918072 $T=13020 4970 0 0 $X=12920 $Y=4720
X214 2 M1_PO_CDNS_7656633918072 $T=13950 4030 0 0 $X=13850 $Y=3780
X215 7 M1_PO_CDNS_7656633918072 $T=14880 3560 0 0 $X=14780 $Y=3310
X216 10 M1_PO_CDNS_7656633918072 $T=15810 3090 0 0 $X=15710 $Y=2840
X217 12 M1_PO_CDNS_7656633918072 $T=17670 6850 0 0 $X=17570 $Y=6600
X218 9 M1_PO_CDNS_7656633918072 $T=18600 6380 0 0 $X=18500 $Y=6130
X219 6 M1_PO_CDNS_7656633918072 $T=19530 5910 0 0 $X=19430 $Y=5660
X220 1 M1_PO_CDNS_7656633918072 $T=20460 5440 0 0 $X=20360 $Y=5190
X221 3 M1_PO_CDNS_7656633918072 $T=21390 4970 0 0 $X=21290 $Y=4720
X222 2 M1_PO_CDNS_7656633918072 $T=22320 4030 0 0 $X=22220 $Y=3780
X223 7 M1_PO_CDNS_7656633918072 $T=23250 3560 0 0 $X=23150 $Y=3310
X224 10 M1_PO_CDNS_7656633918072 $T=24180 3090 0 0 $X=24080 $Y=2840
X225 14 M1_PO_CDNS_7656633918072 $T=25110 2620 0 0 $X=25010 $Y=2370
X226 1 M2_M1_CDNS_7656633918074 $T=80 5580 0 0 $X=0 $Y=5190
X227 16 M2_M1_CDNS_7656633918074 $T=1540 7840 0 0 $X=1460 $Y=7450
X228 6 M2_M1_CDNS_7656633918074 $T=2130 6050 0 0 $X=2050 $Y=5660
X229 16 M2_M1_CDNS_7656633918074 $T=2470 1570 0 0 $X=2390 $Y=1180
X230 17 M2_M1_CDNS_7656633918074 $T=5260 7840 0 0 $X=5180 $Y=7450
X231 17 M2_M1_CDNS_7656633918074 $T=6450 7840 0 0 $X=6370 $Y=7450
X232 17 M2_M1_CDNS_7656633918074 $T=6860 1570 0 0 $X=6780 $Y=1180
X233 9 M2_M1_CDNS_7656633918074 $T=7710 6520 0 0 $X=7630 $Y=6130
X234 17 M2_M1_CDNS_7656633918074 $T=8050 1570 0 0 $X=7970 $Y=1180
X235 18 M2_M1_CDNS_7656633918074 $T=10840 7840 0 0 $X=10760 $Y=7450
X236 18 M2_M1_CDNS_7656633918074 $T=12030 7840 0 0 $X=11950 $Y=7450
X237 18 M2_M1_CDNS_7656633918074 $T=12960 7840 0 0 $X=12880 $Y=7450
X238 18 M2_M1_CDNS_7656633918074 $T=13370 1570 0 0 $X=13290 $Y=1180
X239 18 M2_M1_CDNS_7656633918074 $T=14300 1570 0 0 $X=14220 $Y=1180
X240 18 M2_M1_CDNS_7656633918074 $T=15490 1570 0 0 $X=15410 $Y=1180
X241 12 M2_M1_CDNS_7656633918074 $T=16080 6990 0 0 $X=16000 $Y=6600
X242 19 M2_M1_CDNS_7656633918074 $T=18280 7840 0 0 $X=18200 $Y=7450
X243 19 M2_M1_CDNS_7656633918074 $T=19470 7840 0 0 $X=19390 $Y=7450
X244 19 M2_M1_CDNS_7656633918074 $T=20400 7840 0 0 $X=20320 $Y=7450
X245 19 M2_M1_CDNS_7656633918074 $T=21330 7840 0 0 $X=21250 $Y=7450
X246 19 M2_M1_CDNS_7656633918074 $T=21740 1570 0 0 $X=21660 $Y=1180
X247 19 M2_M1_CDNS_7656633918074 $T=22670 1570 0 0 $X=22590 $Y=1180
X248 19 M2_M1_CDNS_7656633918074 $T=23600 1570 0 0 $X=23520 $Y=1180
X249 19 M2_M1_CDNS_7656633918074 $T=24790 1570 0 0 $X=24710 $Y=1180
X250 16 M7_M6_CDNS_7656633918075 $T=3580 4500 0 0 $X=3360 $Y=4250
X251 17 M7_M6_CDNS_7656633918075 $T=9160 4500 0 0 $X=8940 $Y=4250
X252 18 M7_M6_CDNS_7656633918075 $T=16600 4500 0 0 $X=16380 $Y=4250
X253 19 M7_M6_CDNS_7656633918075 $T=25900 4500 0 0 $X=25680 $Y=4250
X254 16 M6_M5_CDNS_7656633918076 $T=1540 7840 0 0 $X=1460 $Y=7450
X255 16 M6_M5_CDNS_7656633918076 $T=2470 1570 0 0 $X=2390 $Y=1180
X256 17 M6_M5_CDNS_7656633918076 $T=5260 7840 0 0 $X=5180 $Y=7450
X257 17 M6_M5_CDNS_7656633918076 $T=6450 7840 0 0 $X=6370 $Y=7450
X258 17 M6_M5_CDNS_7656633918076 $T=6860 1570 0 0 $X=6780 $Y=1180
X259 17 M6_M5_CDNS_7656633918076 $T=8050 1570 0 0 $X=7970 $Y=1180
X260 18 M6_M5_CDNS_7656633918076 $T=10840 7840 0 0 $X=10760 $Y=7450
X261 18 M6_M5_CDNS_7656633918076 $T=12030 7840 0 0 $X=11950 $Y=7450
X262 18 M6_M5_CDNS_7656633918076 $T=12960 7840 0 0 $X=12880 $Y=7450
X263 18 M6_M5_CDNS_7656633918076 $T=13370 1570 0 0 $X=13290 $Y=1180
X264 18 M6_M5_CDNS_7656633918076 $T=14300 1570 0 0 $X=14220 $Y=1180
X265 18 M6_M5_CDNS_7656633918076 $T=15490 1570 0 0 $X=15410 $Y=1180
X266 19 M6_M5_CDNS_7656633918076 $T=18280 7840 0 0 $X=18200 $Y=7450
X267 19 M6_M5_CDNS_7656633918076 $T=19470 7840 0 0 $X=19390 $Y=7450
X268 19 M6_M5_CDNS_7656633918076 $T=20400 7840 0 0 $X=20320 $Y=7450
X269 19 M6_M5_CDNS_7656633918076 $T=21330 7840 0 0 $X=21250 $Y=7450
X270 19 M6_M5_CDNS_7656633918076 $T=21740 1570 0 0 $X=21660 $Y=1180
X271 19 M6_M5_CDNS_7656633918076 $T=22670 1570 0 0 $X=22590 $Y=1180
X272 19 M6_M5_CDNS_7656633918076 $T=23600 1570 0 0 $X=23520 $Y=1180
X273 19 M6_M5_CDNS_7656633918076 $T=24790 1570 0 0 $X=24710 $Y=1180
X274 1 M6_M5_CDNS_7656633918077 $T=80 5580 0 0 $X=0 $Y=5190
X275 6 M6_M5_CDNS_7656633918077 $T=2130 6050 0 0 $X=2050 $Y=5660
X276 9 M6_M5_CDNS_7656633918077 $T=7710 6520 0 0 $X=7630 $Y=6130
X277 12 M6_M5_CDNS_7656633918077 $T=16080 6990 0 0 $X=16000 $Y=6600
X278 1 M3_M2_CDNS_7656633918078 $T=80 5580 0 0 $X=0 $Y=5190
X279 16 M3_M2_CDNS_7656633918078 $T=1540 7840 0 0 $X=1460 $Y=7450
X280 6 M3_M2_CDNS_7656633918078 $T=2130 6050 0 0 $X=2050 $Y=5660
X281 16 M3_M2_CDNS_7656633918078 $T=2470 1570 0 0 $X=2390 $Y=1180
X282 17 M3_M2_CDNS_7656633918078 $T=5260 7840 0 0 $X=5180 $Y=7450
X283 17 M3_M2_CDNS_7656633918078 $T=6450 7840 0 0 $X=6370 $Y=7450
X284 17 M3_M2_CDNS_7656633918078 $T=6860 1570 0 0 $X=6780 $Y=1180
X285 9 M3_M2_CDNS_7656633918078 $T=7710 6520 0 0 $X=7630 $Y=6130
X286 17 M3_M2_CDNS_7656633918078 $T=8050 1570 0 0 $X=7970 $Y=1180
X287 18 M3_M2_CDNS_7656633918078 $T=10840 7840 0 0 $X=10760 $Y=7450
X288 18 M3_M2_CDNS_7656633918078 $T=12030 7840 0 0 $X=11950 $Y=7450
X289 18 M3_M2_CDNS_7656633918078 $T=12960 7840 0 0 $X=12880 $Y=7450
X290 18 M3_M2_CDNS_7656633918078 $T=13370 1570 0 0 $X=13290 $Y=1180
X291 18 M3_M2_CDNS_7656633918078 $T=14300 1570 0 0 $X=14220 $Y=1180
X292 18 M3_M2_CDNS_7656633918078 $T=15490 1570 0 0 $X=15410 $Y=1180
X293 12 M3_M2_CDNS_7656633918078 $T=16080 6990 0 0 $X=16000 $Y=6600
X294 19 M3_M2_CDNS_7656633918078 $T=18280 7840 0 0 $X=18200 $Y=7450
X295 19 M3_M2_CDNS_7656633918078 $T=19470 7840 0 0 $X=19390 $Y=7450
X296 19 M3_M2_CDNS_7656633918078 $T=20400 7840 0 0 $X=20320 $Y=7450
X297 19 M3_M2_CDNS_7656633918078 $T=21330 7840 0 0 $X=21250 $Y=7450
X298 19 M3_M2_CDNS_7656633918078 $T=21740 1570 0 0 $X=21660 $Y=1180
X299 19 M3_M2_CDNS_7656633918078 $T=22670 1570 0 0 $X=22590 $Y=1180
X300 19 M3_M2_CDNS_7656633918078 $T=23600 1570 0 0 $X=23520 $Y=1180
X301 19 M3_M2_CDNS_7656633918078 $T=24790 1570 0 0 $X=24710 $Y=1180
X302 1 M5_M4_CDNS_7656633918079 $T=80 5580 0 0 $X=0 $Y=5190
X303 16 M5_M4_CDNS_7656633918079 $T=1540 7840 0 0 $X=1460 $Y=7450
X304 6 M5_M4_CDNS_7656633918079 $T=2130 6050 0 0 $X=2050 $Y=5660
X305 16 M5_M4_CDNS_7656633918079 $T=2470 1570 0 0 $X=2390 $Y=1180
X306 17 M5_M4_CDNS_7656633918079 $T=5260 7840 0 0 $X=5180 $Y=7450
X307 17 M5_M4_CDNS_7656633918079 $T=6450 7840 0 0 $X=6370 $Y=7450
X308 17 M5_M4_CDNS_7656633918079 $T=6860 1570 0 0 $X=6780 $Y=1180
X309 9 M5_M4_CDNS_7656633918079 $T=7710 6520 0 0 $X=7630 $Y=6130
X310 17 M5_M4_CDNS_7656633918079 $T=8050 1570 0 0 $X=7970 $Y=1180
X311 18 M5_M4_CDNS_7656633918079 $T=10840 7840 0 0 $X=10760 $Y=7450
X312 18 M5_M4_CDNS_7656633918079 $T=12030 7840 0 0 $X=11950 $Y=7450
X313 18 M5_M4_CDNS_7656633918079 $T=12960 7840 0 0 $X=12880 $Y=7450
X314 18 M5_M4_CDNS_7656633918079 $T=13370 1570 0 0 $X=13290 $Y=1180
X315 18 M5_M4_CDNS_7656633918079 $T=14300 1570 0 0 $X=14220 $Y=1180
X316 18 M5_M4_CDNS_7656633918079 $T=15490 1570 0 0 $X=15410 $Y=1180
X317 12 M5_M4_CDNS_7656633918079 $T=16080 6990 0 0 $X=16000 $Y=6600
X318 19 M5_M4_CDNS_7656633918079 $T=18280 7840 0 0 $X=18200 $Y=7450
X319 19 M5_M4_CDNS_7656633918079 $T=19470 7840 0 0 $X=19390 $Y=7450
X320 19 M5_M4_CDNS_7656633918079 $T=20400 7840 0 0 $X=20320 $Y=7450
X321 19 M5_M4_CDNS_7656633918079 $T=21330 7840 0 0 $X=21250 $Y=7450
X322 19 M5_M4_CDNS_7656633918079 $T=21740 1570 0 0 $X=21660 $Y=1180
X323 19 M5_M4_CDNS_7656633918079 $T=22670 1570 0 0 $X=22590 $Y=1180
X324 19 M5_M4_CDNS_7656633918079 $T=23600 1570 0 0 $X=23520 $Y=1180
X325 19 M5_M4_CDNS_7656633918079 $T=24790 1570 0 0 $X=24710 $Y=1180
X326 4 4 1 16 5 pmos1v_CDNS_7656633918019 $T=1030 8610 1 0 $X=610 $Y=8170
X327 20 4 3 16 5 pmos1v_CDNS_7656633918019 $T=2050 8610 0 180 $X=1540 $Y=8170
X328 22 4 1 17 5 pmos1v_CDNS_7656633918019 $T=5770 8610 0 180 $X=5260 $Y=8170
X329 4 4 18 13 5 pmos1v_CDNS_7656633918019 $T=16840 8610 1 0 $X=16420 $Y=8170
X330 29 4 9 19 5 pmos1v_CDNS_7656633918019 $T=18790 8610 0 180 $X=18280 $Y=8170
X331 28 4 3 19 5 pmos1v_CDNS_7656633918019 $T=21580 8610 0 180 $X=21070 $Y=8170
X332 29 4 10 26 5 pmos1v_CDNS_7656633918019 $T=24370 8610 0 180 $X=23860 $Y=8170
X333 5 5 2 16 nmos1v_CDNS_7656633918020 $T=2980 1040 0 180 $X=2470 $Y=240
X334 5 5 16 8 nmos1v_CDNS_7656633918020 $T=3820 1040 1 0 $X=3400 $Y=240
X335 31 5 1 37 nmos1v_CDNS_7656633918020 $T=5680 1040 1 0 $X=5260 $Y=240
X336 37 5 3 17 nmos1v_CDNS_7656633918020 $T=6610 1040 1 0 $X=6190 $Y=240
X337 5 5 9 34 nmos1v_CDNS_7656633918020 $T=10330 1040 1 0 $X=9910 $Y=240
X338 34 5 6 32 nmos1v_CDNS_7656633918020 $T=11260 1040 1 0 $X=10840 $Y=240
X339 32 5 2 18 nmos1v_CDNS_7656633918020 $T=14050 1040 1 0 $X=13630 $Y=240
X340 5 5 12 35 nmos1v_CDNS_7656633918020 $T=17770 1040 1 0 $X=17350 $Y=240
X341 36 5 6 38 nmos1v_CDNS_7656633918020 $T=19630 1040 1 0 $X=19210 $Y=240
X342 38 5 1 39 nmos1v_CDNS_7656633918020 $T=20560 1040 1 0 $X=20140 $Y=240
X343 39 5 3 19 nmos1v_CDNS_7656633918020 $T=21490 1040 1 0 $X=21070 $Y=240
X344 38 5 2 19 nmos1v_CDNS_7656633918020 $T=22420 1040 1 0 $X=22000 $Y=240
X345 35 5 10 19 nmos1v_CDNS_7656633918020 $T=24280 1040 1 0 $X=23860 $Y=240
X346 5 5 14 19 nmos1v_CDNS_7656633918020 $T=25300 1040 0 180 $X=24790 $Y=240
M0 30 1 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1030 $Y=800 $dt=0
M1 16 3 30 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1960 $Y=800 $dt=0
M2 31 6 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=4750 $Y=800 $dt=0
M3 17 2 31 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=7540 $Y=800 $dt=0
M4 5 7 17 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=8470 $Y=800 $dt=0
M5 11 17 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=9400 $Y=800 $dt=0
M6 33 1 32 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12190 $Y=800 $dt=0
M7 18 3 33 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=13120 $Y=800 $dt=0
M8 18 7 34 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=14980 $Y=800 $dt=0
M9 5 10 18 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=15910 $Y=800 $dt=0
M10 13 18 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=16840 $Y=800 $dt=0
M11 36 9 35 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=18700 $Y=800 $dt=0
M12 19 7 36 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=23350 $Y=800 $dt=0
M13 15 19 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=26140 $Y=800 $dt=0
M14 16 1 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=1030 $Y=8370 $dt=1
M15 20 3 16 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=1960 $Y=8370 $dt=1
M16 4 2 20 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M17 8 16 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M18 17 6 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M19 22 1 17 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=5680 $Y=8370 $dt=1
M20 21 3 17 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M21 22 2 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M22 4 7 22 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M23 11 17 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M24 18 9 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M25 23 6 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M26 24 1 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M27 25 3 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M28 24 2 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M29 23 7 24 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M30 4 10 23 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M31 13 18 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=16840 $Y=8370 $dt=1
M32 19 12 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M33 29 9 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=18700 $Y=8370 $dt=1
M34 26 6 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M35 27 1 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M36 28 3 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=21490 $Y=8370 $dt=1
M37 27 2 28 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M38 26 7 27 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
M39 29 10 26 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=24280 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceFinalAdder                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceFinalAdder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58
** N=164 EP=58 FDC=320
X0 33 M4_M3_CDNS_7656633918010 $T=150 2650 0 0 $X=70 $Y=2400
X1 34 M4_M3_CDNS_7656633918010 $T=5940 2650 0 0 $X=5860 $Y=2400
X2 35 M4_M3_CDNS_7656633918010 $T=16170 2650 0 0 $X=16090 $Y=2400
X3 36 M4_M3_CDNS_7656633918010 $T=21750 2650 0 0 $X=21670 $Y=2400
X4 37 M4_M3_CDNS_7656633918010 $T=26890 2650 0 0 $X=26810 $Y=2400
X5 38 M4_M3_CDNS_7656633918010 $T=32670 2650 0 0 $X=32590 $Y=2400
X6 39 M4_M3_CDNS_7656633918010 $T=40090 2650 0 0 $X=40010 $Y=2400
X7 40 M4_M3_CDNS_7656633918010 $T=48440 2650 0 0 $X=48360 $Y=2400
X8 41 M4_M3_CDNS_7656633918010 $T=53580 2650 0 0 $X=53500 $Y=2400
X9 33 M3_M2_CDNS_7656633918011 $T=150 2650 0 0 $X=70 $Y=2400
X10 34 M3_M2_CDNS_7656633918011 $T=5940 2650 0 0 $X=5860 $Y=2400
X11 35 M3_M2_CDNS_7656633918011 $T=16170 2650 0 0 $X=16090 $Y=2400
X12 36 M3_M2_CDNS_7656633918011 $T=21750 2650 0 0 $X=21670 $Y=2400
X13 37 M3_M2_CDNS_7656633918011 $T=26890 2650 0 0 $X=26810 $Y=2400
X14 38 M3_M2_CDNS_7656633918011 $T=32670 2650 0 0 $X=32590 $Y=2400
X15 39 M3_M2_CDNS_7656633918011 $T=40090 2650 0 0 $X=40010 $Y=2400
X16 40 M3_M2_CDNS_7656633918011 $T=48440 2650 0 0 $X=48360 $Y=2400
X17 41 M3_M2_CDNS_7656633918011 $T=53580 2650 0 0 $X=53500 $Y=2400
X18 1 M2_M1_CDNS_7656633918020 $T=4820 20240 0 0 $X=4740 $Y=20110
X19 9 M2_M1_CDNS_7656633918020 $T=13610 20240 0 0 $X=13530 $Y=20110
X20 12 M2_M1_CDNS_7656633918020 $T=19200 20240 0 0 $X=19120 $Y=20110
X21 17 M2_M1_CDNS_7656633918020 $T=31060 20240 0 0 $X=30980 $Y=20110
X22 18 M2_M1_CDNS_7656633918020 $T=31510 20240 0 0 $X=31430 $Y=20110
X23 21 M2_M1_CDNS_7656633918020 $T=40300 20240 0 0 $X=40220 $Y=20110
X24 24 M2_M1_CDNS_7656633918020 $T=45890 20240 0 0 $X=45810 $Y=20110
X25 29 M2_M1_CDNS_7656633918020 $T=57710 20240 0 0 $X=57630 $Y=20110
X26 42 M3_M2_CDNS_7656633918035 $T=560 3210 0 0 $X=480 $Y=2960
X27 43 M3_M2_CDNS_7656633918035 $T=9840 3210 0 0 $X=9760 $Y=2960
X28 44 M3_M2_CDNS_7656633918035 $T=17280 3210 0 0 $X=17200 $Y=2960
X29 45 M3_M2_CDNS_7656633918035 $T=22860 3210 0 0 $X=22780 $Y=2960
X30 46 M3_M2_CDNS_7656633918035 $T=27230 3210 0 0 $X=27150 $Y=2960
X31 47 M3_M2_CDNS_7656633918035 $T=36530 3210 0 0 $X=36450 $Y=2960
X32 48 M3_M2_CDNS_7656633918035 $T=43970 3210 0 0 $X=43890 $Y=2960
X33 49 M3_M2_CDNS_7656633918035 $T=49550 3210 0 0 $X=49470 $Y=2960
X34 42 M4_M3_CDNS_7656633918036 $T=560 3210 0 0 $X=480 $Y=2960
X35 43 M4_M3_CDNS_7656633918036 $T=9840 3210 0 0 $X=9760 $Y=2960
X36 44 M4_M3_CDNS_7656633918036 $T=17280 3210 0 0 $X=17200 $Y=2960
X37 45 M4_M3_CDNS_7656633918036 $T=22860 3210 0 0 $X=22780 $Y=2960
X38 46 M4_M3_CDNS_7656633918036 $T=27230 3210 0 0 $X=27150 $Y=2960
X39 47 M4_M3_CDNS_7656633918036 $T=36530 3210 0 0 $X=36450 $Y=2960
X40 48 M4_M3_CDNS_7656633918036 $T=43970 3210 0 0 $X=43890 $Y=2960
X41 49 M4_M3_CDNS_7656633918036 $T=49550 3210 0 0 $X=49470 $Y=2960
X42 33 M5_M4_CDNS_7656633918045 $T=150 2650 0 0 $X=70 $Y=2400
X43 34 M5_M4_CDNS_7656633918045 $T=5940 2650 0 0 $X=5860 $Y=2400
X44 35 M5_M4_CDNS_7656633918045 $T=16170 2650 0 0 $X=16090 $Y=2400
X45 36 M5_M4_CDNS_7656633918045 $T=21750 2650 0 0 $X=21670 $Y=2400
X46 37 M5_M4_CDNS_7656633918045 $T=26890 2650 0 0 $X=26810 $Y=2400
X47 38 M5_M4_CDNS_7656633918045 $T=32670 2650 0 0 $X=32590 $Y=2400
X48 39 M5_M4_CDNS_7656633918045 $T=40090 2650 0 0 $X=40010 $Y=2400
X49 40 M5_M4_CDNS_7656633918045 $T=48440 2650 0 0 $X=48360 $Y=2400
X50 41 M5_M4_CDNS_7656633918045 $T=53580 2650 0 0 $X=53500 $Y=2400
X51 33 M6_M5_CDNS_7656633918053 $T=150 2650 0 0 $X=70 $Y=2400
X52 34 M6_M5_CDNS_7656633918053 $T=5940 2650 0 0 $X=5860 $Y=2400
X53 35 M6_M5_CDNS_7656633918053 $T=16170 2650 0 0 $X=16090 $Y=2400
X54 36 M6_M5_CDNS_7656633918053 $T=21750 2650 0 0 $X=21670 $Y=2400
X55 37 M6_M5_CDNS_7656633918053 $T=26890 2650 0 0 $X=26810 $Y=2400
X56 38 M6_M5_CDNS_7656633918053 $T=32670 2650 0 0 $X=32590 $Y=2400
X57 39 M6_M5_CDNS_7656633918053 $T=40090 2650 0 0 $X=40010 $Y=2400
X58 40 M6_M5_CDNS_7656633918053 $T=48440 2650 0 0 $X=48360 $Y=2400
X59 41 M6_M5_CDNS_7656633918053 $T=53580 2650 0 0 $X=53500 $Y=2400
X60 50 M5_M4_CDNS_7656633918057 $T=9340 19910 0 0 $X=9120 $Y=19660
X61 51 M5_M4_CDNS_7656633918057 $T=18130 19910 0 0 $X=17910 $Y=19660
X62 52 M5_M4_CDNS_7656633918057 $T=23720 19910 0 0 $X=23500 $Y=19660
X63 53 M5_M4_CDNS_7656633918057 $T=26500 19910 0 0 $X=26280 $Y=19660
X64 54 M5_M4_CDNS_7656633918057 $T=36030 19910 0 0 $X=35810 $Y=19660
X65 55 M5_M4_CDNS_7656633918057 $T=44820 19910 0 0 $X=44600 $Y=19660
X66 56 M5_M4_CDNS_7656633918057 $T=50410 19910 0 0 $X=50190 $Y=19660
X67 57 M5_M4_CDNS_7656633918057 $T=53190 19910 0 0 $X=52970 $Y=19660
X68 50 M4_M3_CDNS_7656633918058 $T=9340 19910 0 0 $X=9120 $Y=19660
X69 51 M4_M3_CDNS_7656633918058 $T=18130 19910 0 0 $X=17910 $Y=19660
X70 52 M4_M3_CDNS_7656633918058 $T=23720 19910 0 0 $X=23500 $Y=19660
X71 53 M4_M3_CDNS_7656633918058 $T=26500 19910 0 0 $X=26280 $Y=19660
X72 54 M4_M3_CDNS_7656633918058 $T=36030 19910 0 0 $X=35810 $Y=19660
X73 55 M4_M3_CDNS_7656633918058 $T=44820 19910 0 0 $X=44600 $Y=19660
X74 56 M4_M3_CDNS_7656633918058 $T=50410 19910 0 0 $X=50190 $Y=19660
X75 57 M4_M3_CDNS_7656633918058 $T=53190 19910 0 0 $X=52970 $Y=19660
X76 50 M3_M2_CDNS_7656633918059 $T=9340 19910 0 0 $X=9120 $Y=19660
X77 51 M3_M2_CDNS_7656633918059 $T=18130 19910 0 0 $X=17910 $Y=19660
X78 52 M3_M2_CDNS_7656633918059 $T=23720 19910 0 0 $X=23500 $Y=19660
X79 53 M3_M2_CDNS_7656633918059 $T=26500 19910 0 0 $X=26280 $Y=19660
X80 54 M3_M2_CDNS_7656633918059 $T=36030 19910 0 0 $X=35810 $Y=19660
X81 55 M3_M2_CDNS_7656633918059 $T=44820 19910 0 0 $X=44600 $Y=19660
X82 56 M3_M2_CDNS_7656633918059 $T=50410 19910 0 0 $X=50190 $Y=19660
X83 57 M3_M2_CDNS_7656633918059 $T=53190 19910 0 0 $X=52970 $Y=19660
X84 50 M2_M1_CDNS_7656633918060 $T=9340 19910 0 0 $X=9120 $Y=19660
X85 51 M2_M1_CDNS_7656633918060 $T=18130 19910 0 0 $X=17910 $Y=19660
X86 52 M2_M1_CDNS_7656633918060 $T=23720 19910 0 0 $X=23500 $Y=19660
X87 53 M2_M1_CDNS_7656633918060 $T=26500 19910 0 0 $X=26280 $Y=19660
X88 54 M2_M1_CDNS_7656633918060 $T=36030 19910 0 0 $X=35810 $Y=19660
X89 55 M2_M1_CDNS_7656633918060 $T=44820 19910 0 0 $X=44600 $Y=19660
X90 56 M2_M1_CDNS_7656633918060 $T=50410 19910 0 0 $X=50190 $Y=19660
X91 57 M2_M1_CDNS_7656633918060 $T=53190 19910 0 0 $X=52970 $Y=19660
X92 50 M6_M5_CDNS_7656633918061 $T=9340 19910 0 0 $X=9120 $Y=19660
X93 51 M6_M5_CDNS_7656633918061 $T=18130 19910 0 0 $X=17910 $Y=19660
X94 52 M6_M5_CDNS_7656633918061 $T=23720 19910 0 0 $X=23500 $Y=19660
X95 53 M6_M5_CDNS_7656633918061 $T=26500 19910 0 0 $X=26280 $Y=19660
X96 54 M6_M5_CDNS_7656633918061 $T=36030 19910 0 0 $X=35810 $Y=19660
X97 55 M6_M5_CDNS_7656633918061 $T=44820 19910 0 0 $X=44600 $Y=19660
X98 56 M6_M5_CDNS_7656633918061 $T=50410 19910 0 0 $X=50190 $Y=19660
X99 57 M6_M5_CDNS_7656633918061 $T=53190 19910 0 0 $X=52970 $Y=19660
X100 7 1 6 5 50 66 109 AND $T=3670 21910 0 0 $X=4740 $Y=18810
X101 10 9 6 5 51 70 112 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X102 13 12 6 5 52 73 115 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X103 15 17 6 5 53 80 128 AND $T=32210 21910 1 180 $X=26960 $Y=18810
X104 19 18 6 5 54 82 130 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X105 22 21 6 5 55 86 134 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X106 25 24 6 5 56 89 137 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X107 28 29 6 5 57 94 142 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X108 3 6 5 33 2 106 64 XOR $T=530 18810 1 0 $X=530 $Y=14110
X109 42 6 5 4 33 105 63 XOR $T=640 4700 1 0 $X=640 $Y=0
X110 1 6 5 34 7 108 65 XOR $T=4740 18810 1 0 $X=4740 $Y=14110
X111 43 6 5 8 34 107 67 XOR $T=9740 4700 0 180 $X=6020 $Y=0
X112 44 6 5 11 35 111 69 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X113 9 6 5 35 10 110 68 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X114 45 6 5 14 36 114 72 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X115 12 6 5 36 13 113 71 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X116 46 6 5 16 37 116 74 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X117 17 6 5 37 15 127 79 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X118 18 6 5 38 19 129 81 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X119 47 6 5 20 38 131 83 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X120 48 6 5 23 39 133 85 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X121 21 6 5 39 22 132 84 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X122 49 6 5 27 40 136 88 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X123 24 6 5 40 25 135 87 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X124 58 6 5 26 41 138 90 XOR $T=49650 4700 1 0 $X=49650 $Y=0
X125 29 6 5 41 28 141 93 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X126 30 5 58 31 32 6 92 91 139 163
+ 164 140 HAdder $T=62720 6180 1 90 $X=53760 $Y=6980
X127 37 53 46 6 5 36 52 45 35 51
+ 44 34 43 50 42 59 60 61 62 143
+ 145 144 146 147 148 150 151 152 149 95
+ 96 99 100 98 101 102 97 103 104 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X128 41 57 58 6 5 40 56 49 39 55
+ 48 38 47 54 46 75 76 77 78 153
+ 155 154 156 157 158 160 161 162 159 117
+ 118 121 122 120 123 124 119 125 126 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
M0 109 1 66 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5600 $Y=19150 $dt=0
M1 5 7 109 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5810 $Y=19150 $dt=0
M2 50 66 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=8230 $Y=19140 $dt=0
M3 112 9 70 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=19150 $dt=0
M4 5 10 112 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=19150 $dt=0
M5 51 70 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=19140 $dt=0
M6 115 12 73 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=19150 $dt=0
M7 5 13 115 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=19150 $dt=0
M8 52 73 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=19140 $dt=0
M9 5 80 53 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27560 $Y=19140 $dt=0
M10 128 15 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29980 $Y=19150 $dt=0
M11 80 17 128 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30190 $Y=19150 $dt=0
M12 130 18 82 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=19150 $dt=0
M13 5 19 130 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=19150 $dt=0
M14 54 82 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=19140 $dt=0
M15 134 21 86 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=19150 $dt=0
M16 5 22 134 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=19150 $dt=0
M17 55 86 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=19140 $dt=0
M18 137 24 89 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=19150 $dt=0
M19 5 25 137 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=19150 $dt=0
M20 56 89 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=19140 $dt=0
M21 5 94 57 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=19140 $dt=0
M22 142 28 5 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=19150 $dt=0
M23 94 29 142 5 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=19150 $dt=0
M24 6 62 42 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M25 106 3 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=950 $Y=14910 $dt=1
M26 105 42 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=115.144 scb=0.0588049 scc=0.0138331 $X=1060 $Y=800 $dt=1
M27 149 50 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M28 33 2 3 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=1880 $Y=14910 $dt=1
M29 4 33 42 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.854 scb=0.0354545 scc=0.011187 $X=1990 $Y=800 $dt=1
M30 106 64 33 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=2810 $Y=14910 $dt=1
M31 105 63 4 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=2920 $Y=800 $dt=1
M32 6 2 64 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=3740 $Y=14910 $dt=1
M33 6 33 63 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=3850 $Y=800 $dt=1
M34 108 1 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=14910 $dt=1
M35 66 1 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=20590 $dt=1
M36 6 7 66 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=20590 $dt=1
M37 34 7 1 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=14910 $dt=1
M38 67 34 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=6440 $Y=800 $dt=1
M39 108 65 34 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=14910 $dt=1
M40 8 67 107 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=7370 $Y=800 $dt=1
M41 6 7 65 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=14910 $dt=1
M42 50 66 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=8230 $Y=20400 $dt=1
M43 43 34 8 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=8300 $Y=800 $dt=1
M44 6 43 107 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=9230 $Y=800 $dt=1
M45 69 35 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=13880 $Y=800 $dt=1
M46 110 9 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M47 70 9 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=20590 $dt=1
M48 6 10 70 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=20590 $dt=1
M49 11 69 111 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=14810 $Y=800 $dt=1
M50 35 10 9 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M51 44 35 11 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=15740 $Y=800 $dt=1
M52 110 68 35 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M53 6 44 111 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=16670 $Y=800 $dt=1
M54 6 10 68 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M55 51 70 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17020 $Y=20400 $dt=1
M56 72 36 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=19460 $Y=800 $dt=1
M57 113 12 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M58 73 12 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=20590 $dt=1
M59 14 72 114 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=20390 $Y=800 $dt=1
M60 6 13 73 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=20590 $dt=1
M61 36 13 12 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M62 45 36 14 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=21320 $Y=800 $dt=1
M63 113 71 36 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M64 6 45 114 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=22250 $Y=800 $dt=1
M65 6 13 71 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M66 52 73 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22610 $Y=20400 $dt=1
M67 74 37 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=23510 $Y=800 $dt=1
M68 16 74 116 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=24440 $Y=800 $dt=1
M69 46 37 16 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=25370 $Y=800 $dt=1
M70 6 46 116 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=26300 $Y=800 $dt=1
M71 6 78 46 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M72 6 80 53 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27560 $Y=20400 $dt=1
M73 79 15 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M74 159 54 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M75 37 79 127 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M76 17 15 37 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M77 80 15 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29780 $Y=20590 $dt=1
M78 6 17 80 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30190 $Y=20590 $dt=1
M79 6 17 127 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M80 129 18 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M81 82 18 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=20590 $dt=1
M82 6 19 82 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=20590 $dt=1
M83 38 19 18 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M84 83 38 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=33170 $Y=800 $dt=1
M85 129 81 38 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M86 20 83 131 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=34100 $Y=800 $dt=1
M87 6 19 81 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M88 54 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=34920 $Y=20400 $dt=1
M89 47 38 20 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35030 $Y=800 $dt=1
M90 6 47 131 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35960 $Y=800 $dt=1
M91 85 39 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=40590 $Y=800 $dt=1
M92 132 21 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M93 86 21 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=20590 $dt=1
M94 6 22 86 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=20590 $dt=1
M95 23 85 133 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=41520 $Y=800 $dt=1
M96 39 22 21 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M97 48 39 23 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=42450 $Y=800 $dt=1
M98 132 84 39 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M99 6 48 133 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=43380 $Y=800 $dt=1
M100 6 22 84 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M101 55 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=43710 $Y=20400 $dt=1
M102 88 40 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=46150 $Y=800 $dt=1
M103 135 24 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M104 89 24 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=20590 $dt=1
M105 27 88 136 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=47080 $Y=800 $dt=1
M106 6 25 89 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=20590 $dt=1
M107 40 25 24 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M108 49 40 27 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48010 $Y=800 $dt=1
M109 135 87 40 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M110 6 49 136 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48940 $Y=800 $dt=1
M111 6 25 87 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M112 56 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=49300 $Y=20400 $dt=1
M113 138 58 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=50070 $Y=800 $dt=1
M114 26 41 58 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51000 $Y=800 $dt=1
M115 138 90 26 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51930 $Y=800 $dt=1
M116 6 41 90 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=52860 $Y=800 $dt=1
M117 6 94 57 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=54210 $Y=20400 $dt=1
M118 93 28 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M119 41 93 141 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M120 164 92 58 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=55830 $Y=11700 $dt=1
M121 6 91 164 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56040 $Y=11700 $dt=1
M122 29 28 41 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M123 94 28 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=20590 $dt=1
M124 6 29 94 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=20590 $dt=1
M125 6 91 163 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56970 $Y=11700 $dt=1
M126 6 29 141 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M127 163 92 6 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57380 $Y=11700 $dt=1
M128 30 32 163 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57790 $Y=11700 $dt=1
M129 163 31 30 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=58200 $Y=11700 $dt=1
M130 6 31 91 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=59130 $Y=11700 $dt=1
M131 6 32 92 6 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=60060 $Y=11700 $dt=1
.ends WallaceFinalAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_7656633918080                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_7656633918080 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_7656633918080

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918021                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918021 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656633918021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918022                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918022 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656633918022

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918023                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918023 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_7656633918023

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656633918024                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656633918024 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_7656633918024

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918025                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918025 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.6986 scb=0.0347897 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656633918025

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918026                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918026 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656633918026

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656633918027                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656633918027 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656633918027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAdder 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=10
X0 8 M2_M1_CDNS_7656633918020 $T=2700 5110 0 90 $X=2570 $Y=5030
X1 9 M2_M1_CDNS_7656633918020 $T=3060 2950 0 90 $X=2930 $Y=2870
X2 9 M2_M1_CDNS_7656633918020 $T=3060 5520 0 90 $X=2930 $Y=5440
X3 5 M2_M1_CDNS_7656633918020 $T=3450 7370 0 90 $X=3320 $Y=7290
X4 3 M2_M1_CDNS_7656633918020 $T=3450 8190 0 90 $X=3320 $Y=8110
X5 5 M2_M1_CDNS_7656633918020 $T=3460 3880 0 90 $X=3330 $Y=3800
X6 3 M2_M1_CDNS_7656633918020 $T=4250 4700 0 90 $X=4120 $Y=4620
X7 10 M2_M1_CDNS_7656633918020 $T=4700 5110 0 90 $X=4570 $Y=5030
X8 10 M2_M1_CDNS_7656633918020 $T=4740 5820 0 90 $X=4610 $Y=5740
X9 8 M2_M1_CDNS_7656633918020 $T=5140 5990 0 90 $X=5010 $Y=5910
X10 8 M2_M1_CDNS_7656633918025 $T=5020 6720 0 90 $X=4890 $Y=6590
X11 10 M1_PO_CDNS_7656633918062 $T=1550 6040 0 90 $X=1430 $Y=5940
X12 5 M1_PO_CDNS_7656633918062 $T=3090 2650 0 90 $X=2970 $Y=2550
X13 5 M1_PO_CDNS_7656633918062 $T=3090 3820 0 90 $X=2970 $Y=3720
X14 5 M1_PO_CDNS_7656633918062 $T=3090 4360 0 90 $X=2970 $Y=4260
X15 6 M1_PO_CDNS_7656633918062 $T=3145 6870 0 90 $X=3025 $Y=6770
X16 9 M1_PO_CDNS_7656633918062 $T=3720 5020 0 90 $X=3600 $Y=4920
X17 8 M1_PO_CDNS_7656633918063 $T=2700 7470 0 90 $X=2450 $Y=7370
X18 6 M1_PO_CDNS_7656633918063 $T=3820 6180 0 90 $X=3570 $Y=6080
X19 3 M1_PO_CDNS_7656633918063 $T=4200 5220 0 90 $X=3950 $Y=5120
X20 3 M1_PO_CDNS_7656633918063 $T=4250 4170 0 90 $X=4000 $Y=4070
X21 10 M1_PO_CDNS_7656633918063 $T=4650 8090 0 90 $X=4400 $Y=7990
X22 8 M1_PO_CDNS_7656633918063 $T=5020 6720 0 90 $X=4770 $Y=6620
X23 8 M2_M1_CDNS_7656633918064 $T=2700 7470 0 90 $X=2450 $Y=7390
X24 6 M2_M1_CDNS_7656633918064 $T=3820 6180 0 90 $X=3570 $Y=6100
X25 3 M2_M1_CDNS_7656633918064 $T=4200 5220 0 90 $X=3950 $Y=5140
X26 3 M2_M1_CDNS_7656633918064 $T=4250 4170 0 90 $X=4000 $Y=4090
X27 10 M2_M1_CDNS_7656633918064 $T=4650 8090 0 90 $X=4400 $Y=8010
X28 9 3 8 1 nmos1v_CDNS_7656633918014 $T=2220 5270 0 90 $X=1780 $Y=5030
X29 10 6 2 1 nmos1v_CDNS_7656633918014 $T=2220 6290 1 270 $X=1780 $Y=5780
X30 3 10 4 1 nmos1v_CDNS_7656633918014 $T=2220 7950 0 90 $X=1780 $Y=7710
X31 5 3 8 1 7 pmos1v_CDNS_7656633918018 $T=5670 4040 0 90 $X=5230 $Y=3620
X32 9 3 10 1 7 pmos1v_CDNS_7656633918018 $T=5670 5360 1 270 $X=5230 $Y=5030
X33 5 8 4 1 7 pmos1v_CDNS_7656633918018 $T=5670 7540 0 90 $X=5230 $Y=7120
X34 7 7 5 9 1 pmos1v_CDNS_7656633918019 $T=5670 3200 1 270 $X=5230 $Y=2690
X35 1 1 5 9 nmos1v_CDNS_7656633918020 $T=2220 3200 1 270 $X=1420 $Y=2690
X36 6 M2_M1_CDNS_7656633918080 $T=3820 2110 0 90 $X=3740 $Y=1860
X37 3 M2_M1_CDNS_7656633918080 $T=4260 2110 0 90 $X=4180 $Y=1860
X38 5 3 10 1 nmos1v_CDNS_7656633918021 $T=2220 4450 0 90 $X=1780 $Y=4210
X39 10 5 3 1 nmos1v_CDNS_7656633918022 $T=2220 4130 1 270 $X=1780 $Y=3620
X40 2 6 10 1 nmos1v_CDNS_7656633918022 $T=2220 6610 0 90 $X=1780 $Y=6250
X41 4 6 8 1 nmos1v_CDNS_7656633918022 $T=2220 7630 1 270 $X=1780 $Y=7120
X42 6 8 2 1 7 pmos1v_CDNS_7656633918023 $T=5670 6700 1 270 $X=5230 $Y=6250
X43 6 10 4 1 7 pmos1v_CDNS_7656633918023 $T=5670 8040 1 270 $X=5230 $Y=7590
X44 8 3 9 1 nmos1v_CDNS_7656633918024 $T=2220 4950 1 270 $X=1780 $Y=4500
X45 8 5 3 1 7 pmos1v_CDNS_7656633918025 $T=5670 4540 1 270 $X=5230 $Y=4090
X46 3 10 9 1 7 pmos1v_CDNS_7656633918026 $T=5670 4860 0 90 $X=5230 $Y=4500
X47 8 6 2 1 7 pmos1v_CDNS_7656633918027 $T=5670 6200 0 90 $X=5230 $Y=5780
M0 4 8 6 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1980 $Y=7540 $dt=0
M1 7 5 9 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5430 $Y=3110 $dt=1
M2 8 3 5 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5430 $Y=4040 $dt=1
M3 9 3 10 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5430 $Y=5270 $dt=1
M4 6 8 2 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=95.6709 scb=0.0347795 scc=0.0111862 $X=5430 $Y=6610 $dt=1
M5 4 8 5 7 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=99.6807 scb=0.0402027 scc=0.0112574 $X=5430 $Y=7540 $dt=1
.ends FAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y1 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=0
X0 1 M2_M1_CDNS_7656633918028 $T=80 250 0 0 $X=0 $Y=0
X1 2 M2_M1_CDNS_7656633918028 $T=480 250 0 0 $X=400 $Y=0
X2 3 M2_M1_CDNS_7656633918028 $T=880 250 0 0 $X=800 $Y=0
X3 4 M2_M1_CDNS_7656633918028 $T=1280 250 0 0 $X=1200 $Y=0
X4 5 M2_M1_CDNS_7656633918028 $T=1680 250 0 0 $X=1600 $Y=0
X5 6 M2_M1_CDNS_7656633918028 $T=2080 250 0 0 $X=2000 $Y=0
X6 7 M2_M1_CDNS_7656633918028 $T=2480 250 0 0 $X=2400 $Y=0
X7 8 M2_M1_CDNS_7656633918028 $T=2880 250 0 0 $X=2800 $Y=0
.ends MASCO__Y1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__Y2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__Y2 1 2 3 4 5 6 7 8
** N=8 EP=8 FDC=0
X0 1 M3_M2_CDNS_7656633918027 $T=80 250 0 0 $X=0 $Y=0
X1 2 M3_M2_CDNS_7656633918027 $T=480 250 0 0 $X=400 $Y=0
X2 3 M3_M2_CDNS_7656633918027 $T=880 250 0 0 $X=800 $Y=0
X3 4 M3_M2_CDNS_7656633918027 $T=1280 250 0 0 $X=1200 $Y=0
X4 5 M3_M2_CDNS_7656633918027 $T=1680 250 0 0 $X=1600 $Y=0
X5 6 M3_M2_CDNS_7656633918027 $T=2080 250 0 0 $X=2000 $Y=0
X6 7 M3_M2_CDNS_7656633918027 $T=2480 250 0 0 $X=2400 $Y=0
X7 8 M3_M2_CDNS_7656633918027 $T=2880 250 0 0 $X=2800 $Y=0
.ends MASCO__Y2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceMultiplier                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceMultiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82
** N=210 EP=82 FDC=384
X0 2 M2_M1_CDNS_7656633918020 $T=2220 31930 0 0 $X=2140 $Y=31800
X1 3 M2_M1_CDNS_7656633918020 $T=2220 35820 0 0 $X=2140 $Y=35690
X2 4 M2_M1_CDNS_7656633918020 $T=2220 36470 0 0 $X=2140 $Y=36340
X3 5 M2_M1_CDNS_7656633918020 $T=2220 40360 0 0 $X=2140 $Y=40230
X4 6 M2_M1_CDNS_7656633918020 $T=2220 41010 0 0 $X=2140 $Y=40880
X5 7 M2_M1_CDNS_7656633918020 $T=2220 44900 0 0 $X=2140 $Y=44770
X6 8 M2_M1_CDNS_7656633918020 $T=2220 45540 0 0 $X=2140 $Y=45410
X7 9 M2_M1_CDNS_7656633918020 $T=2220 49430 0 0 $X=2140 $Y=49300
X8 2 M2_M1_CDNS_7656633918020 $T=3380 32500 0 0 $X=3300 $Y=32370
X9 3 M2_M1_CDNS_7656633918020 $T=3380 35240 0 0 $X=3300 $Y=35110
X10 4 M2_M1_CDNS_7656633918020 $T=3380 37040 0 0 $X=3300 $Y=36910
X11 5 M2_M1_CDNS_7656633918020 $T=3380 39780 0 0 $X=3300 $Y=39650
X12 6 M2_M1_CDNS_7656633918020 $T=3380 41580 0 0 $X=3300 $Y=41450
X13 7 M2_M1_CDNS_7656633918020 $T=3380 44320 0 0 $X=3300 $Y=44190
X14 8 M2_M1_CDNS_7656633918020 $T=3380 46120 0 0 $X=3300 $Y=45990
X15 9 M2_M1_CDNS_7656633918020 $T=3380 48860 0 0 $X=3300 $Y=48730
X16 2 M2_M1_CDNS_7656633918020 $T=8590 32500 0 0 $X=8510 $Y=32370
X17 3 M2_M1_CDNS_7656633918020 $T=8590 35240 0 0 $X=8510 $Y=35110
X18 4 M2_M1_CDNS_7656633918020 $T=8590 37040 0 0 $X=8510 $Y=36910
X19 5 M2_M1_CDNS_7656633918020 $T=8590 39780 0 0 $X=8510 $Y=39650
X20 6 M2_M1_CDNS_7656633918020 $T=8590 41580 0 0 $X=8510 $Y=41450
X21 7 M2_M1_CDNS_7656633918020 $T=8590 44320 0 0 $X=8510 $Y=44190
X22 8 M2_M1_CDNS_7656633918020 $T=8590 46120 0 0 $X=8510 $Y=45990
X23 9 M2_M1_CDNS_7656633918020 $T=8590 48860 0 0 $X=8510 $Y=48730
X24 2 M2_M1_CDNS_7656633918020 $T=13610 32500 0 0 $X=13530 $Y=32370
X25 3 M2_M1_CDNS_7656633918020 $T=13610 35240 0 0 $X=13530 $Y=35110
X26 4 M2_M1_CDNS_7656633918020 $T=13610 37040 0 0 $X=13530 $Y=36910
X27 5 M2_M1_CDNS_7656633918020 $T=13610 39780 0 0 $X=13530 $Y=39650
X28 6 M2_M1_CDNS_7656633918020 $T=13610 41580 0 0 $X=13530 $Y=41450
X29 7 M2_M1_CDNS_7656633918020 $T=13610 44320 0 0 $X=13530 $Y=44190
X30 8 M2_M1_CDNS_7656633918020 $T=13610 46120 0 0 $X=13530 $Y=45990
X31 9 M2_M1_CDNS_7656633918020 $T=13610 48860 0 0 $X=13530 $Y=48730
X32 2 M2_M1_CDNS_7656633918020 $T=18740 32500 0 0 $X=18660 $Y=32370
X33 3 M2_M1_CDNS_7656633918020 $T=18740 35240 0 0 $X=18660 $Y=35110
X34 4 M2_M1_CDNS_7656633918020 $T=18740 37040 0 0 $X=18660 $Y=36910
X35 5 M2_M1_CDNS_7656633918020 $T=18740 39780 0 0 $X=18660 $Y=39650
X36 6 M2_M1_CDNS_7656633918020 $T=18740 41580 0 0 $X=18660 $Y=41450
X37 7 M2_M1_CDNS_7656633918020 $T=18740 44320 0 0 $X=18660 $Y=44190
X38 8 M2_M1_CDNS_7656633918020 $T=18740 46120 0 0 $X=18660 $Y=45990
X39 9 M2_M1_CDNS_7656633918020 $T=18740 48860 0 0 $X=18660 $Y=48730
X40 2 M2_M1_CDNS_7656633918020 $T=23810 32500 0 0 $X=23730 $Y=32370
X41 3 M2_M1_CDNS_7656633918020 $T=23810 35240 0 0 $X=23730 $Y=35110
X42 4 M2_M1_CDNS_7656633918020 $T=23810 37040 0 0 $X=23730 $Y=36910
X43 5 M2_M1_CDNS_7656633918020 $T=23810 39780 0 0 $X=23730 $Y=39650
X44 6 M2_M1_CDNS_7656633918020 $T=23810 41580 0 0 $X=23730 $Y=41450
X45 7 M2_M1_CDNS_7656633918020 $T=23810 44320 0 0 $X=23730 $Y=44190
X46 8 M2_M1_CDNS_7656633918020 $T=23810 46120 0 0 $X=23730 $Y=45990
X47 9 M2_M1_CDNS_7656633918020 $T=23810 48860 0 0 $X=23730 $Y=48730
X48 2 M2_M1_CDNS_7656633918020 $T=28690 32500 0 0 $X=28610 $Y=32370
X49 3 M2_M1_CDNS_7656633918020 $T=28690 35240 0 0 $X=28610 $Y=35110
X50 4 M2_M1_CDNS_7656633918020 $T=28690 37040 0 0 $X=28610 $Y=36910
X51 5 M2_M1_CDNS_7656633918020 $T=28690 39780 0 0 $X=28610 $Y=39650
X52 6 M2_M1_CDNS_7656633918020 $T=28690 41580 0 0 $X=28610 $Y=41450
X53 7 M2_M1_CDNS_7656633918020 $T=28690 44320 0 0 $X=28610 $Y=44190
X54 8 M2_M1_CDNS_7656633918020 $T=28690 46120 0 0 $X=28610 $Y=45990
X55 9 M2_M1_CDNS_7656633918020 $T=28690 48860 0 0 $X=28610 $Y=48730
X56 2 M2_M1_CDNS_7656633918020 $T=33890 32500 0 0 $X=33810 $Y=32370
X57 3 M2_M1_CDNS_7656633918020 $T=33890 35240 0 0 $X=33810 $Y=35110
X58 4 M2_M1_CDNS_7656633918020 $T=33890 37040 0 0 $X=33810 $Y=36910
X59 5 M2_M1_CDNS_7656633918020 $T=33890 39780 0 0 $X=33810 $Y=39650
X60 6 M2_M1_CDNS_7656633918020 $T=33890 41580 0 0 $X=33810 $Y=41450
X61 7 M2_M1_CDNS_7656633918020 $T=33890 44320 0 0 $X=33810 $Y=44190
X62 8 M2_M1_CDNS_7656633918020 $T=33890 46120 0 0 $X=33810 $Y=45990
X63 9 M2_M1_CDNS_7656633918020 $T=33890 48860 0 0 $X=33810 $Y=48730
X64 2 M2_M1_CDNS_7656633918020 $T=38920 32500 0 0 $X=38840 $Y=32370
X65 3 M2_M1_CDNS_7656633918020 $T=38920 35240 0 0 $X=38840 $Y=35110
X66 4 M2_M1_CDNS_7656633918020 $T=38920 37040 0 0 $X=38840 $Y=36910
X67 5 M2_M1_CDNS_7656633918020 $T=38920 39780 0 0 $X=38840 $Y=39650
X68 6 M2_M1_CDNS_7656633918020 $T=38920 41580 0 0 $X=38840 $Y=41450
X69 7 M2_M1_CDNS_7656633918020 $T=38920 44320 0 0 $X=38840 $Y=44190
X70 8 M2_M1_CDNS_7656633918020 $T=38920 46120 0 0 $X=38840 $Y=45990
X71 9 M2_M1_CDNS_7656633918020 $T=38920 48860 0 0 $X=38840 $Y=48730
X72 1 M3_M2_CDNS_7656633918027 $T=3380 31230 0 0 $X=3300 $Y=30980
X73 1 M3_M2_CDNS_7656633918027 $T=3380 33140 0 0 $X=3300 $Y=32890
X74 1 M3_M2_CDNS_7656633918027 $T=3380 34600 0 0 $X=3300 $Y=34350
X75 1 M3_M2_CDNS_7656633918027 $T=3380 37680 0 0 $X=3300 $Y=37430
X76 1 M3_M2_CDNS_7656633918027 $T=3380 39140 0 0 $X=3300 $Y=38890
X77 1 M3_M2_CDNS_7656633918027 $T=3380 42220 0 0 $X=3300 $Y=41970
X78 1 M3_M2_CDNS_7656633918027 $T=3380 43680 0 0 $X=3300 $Y=43430
X79 1 M3_M2_CDNS_7656633918027 $T=3380 46750 0 0 $X=3300 $Y=46500
X80 1 M3_M2_CDNS_7656633918027 $T=3380 48210 0 0 $X=3300 $Y=47960
X81 18 M3_M2_CDNS_7656633918027 $T=8570 31230 0 0 $X=8490 $Y=30980
X82 18 M3_M2_CDNS_7656633918027 $T=8570 33140 0 0 $X=8490 $Y=32890
X83 18 M3_M2_CDNS_7656633918027 $T=8570 34600 0 0 $X=8490 $Y=34350
X84 18 M3_M2_CDNS_7656633918027 $T=8570 37680 0 0 $X=8490 $Y=37430
X85 18 M3_M2_CDNS_7656633918027 $T=8570 39140 0 0 $X=8490 $Y=38890
X86 18 M3_M2_CDNS_7656633918027 $T=8570 42220 0 0 $X=8490 $Y=41970
X87 18 M3_M2_CDNS_7656633918027 $T=8570 43680 0 0 $X=8490 $Y=43430
X88 18 M3_M2_CDNS_7656633918027 $T=8570 46750 0 0 $X=8490 $Y=46500
X89 18 M3_M2_CDNS_7656633918027 $T=8570 48210 0 0 $X=8490 $Y=47960
X90 26 M3_M2_CDNS_7656633918027 $T=13600 31060 0 0 $X=13520 $Y=30810
X91 26 M3_M2_CDNS_7656633918027 $T=13600 33140 0 0 $X=13520 $Y=32890
X92 26 M3_M2_CDNS_7656633918027 $T=13600 34600 0 0 $X=13520 $Y=34350
X93 26 M3_M2_CDNS_7656633918027 $T=13600 37680 0 0 $X=13520 $Y=37430
X94 26 M3_M2_CDNS_7656633918027 $T=13600 39140 0 0 $X=13520 $Y=38890
X95 26 M3_M2_CDNS_7656633918027 $T=13600 42220 0 0 $X=13520 $Y=41970
X96 26 M3_M2_CDNS_7656633918027 $T=13600 43680 0 0 $X=13520 $Y=43430
X97 26 M3_M2_CDNS_7656633918027 $T=13600 46750 0 0 $X=13520 $Y=46500
X98 26 M3_M2_CDNS_7656633918027 $T=13600 48210 0 0 $X=13520 $Y=47960
X99 35 M3_M2_CDNS_7656633918027 $T=18750 31230 0 0 $X=18670 $Y=30980
X100 35 M3_M2_CDNS_7656633918027 $T=18750 33140 0 0 $X=18670 $Y=32890
X101 35 M3_M2_CDNS_7656633918027 $T=18750 34600 0 0 $X=18670 $Y=34350
X102 35 M3_M2_CDNS_7656633918027 $T=18750 37680 0 0 $X=18670 $Y=37430
X103 35 M3_M2_CDNS_7656633918027 $T=18750 39140 0 0 $X=18670 $Y=38890
X104 35 M3_M2_CDNS_7656633918027 $T=18750 42220 0 0 $X=18670 $Y=41970
X105 35 M3_M2_CDNS_7656633918027 $T=18750 43680 0 0 $X=18670 $Y=43430
X106 35 M3_M2_CDNS_7656633918027 $T=18750 46750 0 0 $X=18670 $Y=46500
X107 35 M3_M2_CDNS_7656633918027 $T=18750 48210 0 0 $X=18670 $Y=47960
X108 44 M3_M2_CDNS_7656633918027 $T=23840 31230 0 0 $X=23760 $Y=30980
X109 44 M3_M2_CDNS_7656633918027 $T=23840 33140 0 0 $X=23760 $Y=32890
X110 44 M3_M2_CDNS_7656633918027 $T=23840 34600 0 0 $X=23760 $Y=34350
X111 44 M3_M2_CDNS_7656633918027 $T=23840 37680 0 0 $X=23760 $Y=37430
X112 44 M3_M2_CDNS_7656633918027 $T=23840 39140 0 0 $X=23760 $Y=38890
X113 44 M3_M2_CDNS_7656633918027 $T=23840 42220 0 0 $X=23760 $Y=41970
X114 44 M3_M2_CDNS_7656633918027 $T=23840 43680 0 0 $X=23760 $Y=43430
X115 44 M3_M2_CDNS_7656633918027 $T=23840 46750 0 0 $X=23760 $Y=46500
X116 44 M3_M2_CDNS_7656633918027 $T=23840 48210 0 0 $X=23760 $Y=47960
X117 53 M3_M2_CDNS_7656633918027 $T=28730 31230 0 0 $X=28650 $Y=30980
X118 53 M3_M2_CDNS_7656633918027 $T=28730 33140 0 0 $X=28650 $Y=32890
X119 53 M3_M2_CDNS_7656633918027 $T=28730 34600 0 0 $X=28650 $Y=34350
X120 53 M3_M2_CDNS_7656633918027 $T=28730 37680 0 0 $X=28650 $Y=37430
X121 53 M3_M2_CDNS_7656633918027 $T=28730 39140 0 0 $X=28650 $Y=38890
X122 53 M3_M2_CDNS_7656633918027 $T=28730 42220 0 0 $X=28650 $Y=41970
X123 53 M3_M2_CDNS_7656633918027 $T=28730 43680 0 0 $X=28650 $Y=43430
X124 53 M3_M2_CDNS_7656633918027 $T=28730 46750 0 0 $X=28650 $Y=46500
X125 53 M3_M2_CDNS_7656633918027 $T=28730 48210 0 0 $X=28650 $Y=47960
X126 62 M3_M2_CDNS_7656633918027 $T=33970 31230 0 0 $X=33890 $Y=30980
X127 62 M3_M2_CDNS_7656633918027 $T=33970 33140 0 0 $X=33890 $Y=32890
X128 62 M3_M2_CDNS_7656633918027 $T=33970 34600 0 0 $X=33890 $Y=34350
X129 62 M3_M2_CDNS_7656633918027 $T=33970 37680 0 0 $X=33890 $Y=37430
X130 62 M3_M2_CDNS_7656633918027 $T=33970 39140 0 0 $X=33890 $Y=38890
X131 62 M3_M2_CDNS_7656633918027 $T=33970 42220 0 0 $X=33890 $Y=41970
X132 62 M3_M2_CDNS_7656633918027 $T=33970 43680 0 0 $X=33890 $Y=43430
X133 62 M3_M2_CDNS_7656633918027 $T=33970 46750 0 0 $X=33890 $Y=46500
X134 62 M3_M2_CDNS_7656633918027 $T=33970 48210 0 0 $X=33890 $Y=47960
X135 71 M3_M2_CDNS_7656633918027 $T=39020 31230 0 0 $X=38940 $Y=30980
X136 71 M3_M2_CDNS_7656633918027 $T=39020 33140 0 0 $X=38940 $Y=32890
X137 71 M3_M2_CDNS_7656633918027 $T=39020 34600 0 0 $X=38940 $Y=34350
X138 71 M3_M2_CDNS_7656633918027 $T=39020 37680 0 0 $X=38940 $Y=37430
X139 71 M3_M2_CDNS_7656633918027 $T=39020 39140 0 0 $X=38940 $Y=38890
X140 71 M3_M2_CDNS_7656633918027 $T=39020 42220 0 0 $X=38940 $Y=41970
X141 71 M3_M2_CDNS_7656633918027 $T=39020 43680 0 0 $X=38940 $Y=43430
X142 71 M3_M2_CDNS_7656633918027 $T=39020 46750 0 0 $X=38940 $Y=46500
X143 71 M3_M2_CDNS_7656633918027 $T=39020 48210 0 0 $X=38940 $Y=47960
X144 1 M2_M1_CDNS_7656633918028 $T=3380 31230 0 0 $X=3300 $Y=30980
X145 1 M2_M1_CDNS_7656633918028 $T=3380 33140 0 0 $X=3300 $Y=32890
X146 1 M2_M1_CDNS_7656633918028 $T=3380 34600 0 0 $X=3300 $Y=34350
X147 1 M2_M1_CDNS_7656633918028 $T=3380 37680 0 0 $X=3300 $Y=37430
X148 1 M2_M1_CDNS_7656633918028 $T=3380 39140 0 0 $X=3300 $Y=38890
X149 1 M2_M1_CDNS_7656633918028 $T=3380 42220 0 0 $X=3300 $Y=41970
X150 1 M2_M1_CDNS_7656633918028 $T=3380 43680 0 0 $X=3300 $Y=43430
X151 1 M2_M1_CDNS_7656633918028 $T=3380 46750 0 0 $X=3300 $Y=46500
X152 1 M2_M1_CDNS_7656633918028 $T=3380 48210 0 0 $X=3300 $Y=47960
X153 18 M2_M1_CDNS_7656633918028 $T=8570 31230 0 0 $X=8490 $Y=30980
X154 18 M2_M1_CDNS_7656633918028 $T=8570 33140 0 0 $X=8490 $Y=32890
X155 18 M2_M1_CDNS_7656633918028 $T=8570 34600 0 0 $X=8490 $Y=34350
X156 18 M2_M1_CDNS_7656633918028 $T=8570 37680 0 0 $X=8490 $Y=37430
X157 18 M2_M1_CDNS_7656633918028 $T=8570 39140 0 0 $X=8490 $Y=38890
X158 18 M2_M1_CDNS_7656633918028 $T=8570 42220 0 0 $X=8490 $Y=41970
X159 18 M2_M1_CDNS_7656633918028 $T=8570 43680 0 0 $X=8490 $Y=43430
X160 18 M2_M1_CDNS_7656633918028 $T=8570 46750 0 0 $X=8490 $Y=46500
X161 18 M2_M1_CDNS_7656633918028 $T=8570 48210 0 0 $X=8490 $Y=47960
X162 26 M2_M1_CDNS_7656633918028 $T=13600 31060 0 0 $X=13520 $Y=30810
X163 26 M2_M1_CDNS_7656633918028 $T=13600 33140 0 0 $X=13520 $Y=32890
X164 26 M2_M1_CDNS_7656633918028 $T=13600 34600 0 0 $X=13520 $Y=34350
X165 26 M2_M1_CDNS_7656633918028 $T=13600 37680 0 0 $X=13520 $Y=37430
X166 26 M2_M1_CDNS_7656633918028 $T=13600 39140 0 0 $X=13520 $Y=38890
X167 26 M2_M1_CDNS_7656633918028 $T=13600 42220 0 0 $X=13520 $Y=41970
X168 26 M2_M1_CDNS_7656633918028 $T=13600 43680 0 0 $X=13520 $Y=43430
X169 26 M2_M1_CDNS_7656633918028 $T=13600 46750 0 0 $X=13520 $Y=46500
X170 26 M2_M1_CDNS_7656633918028 $T=13600 48210 0 0 $X=13520 $Y=47960
X171 35 M2_M1_CDNS_7656633918028 $T=18750 31230 0 0 $X=18670 $Y=30980
X172 35 M2_M1_CDNS_7656633918028 $T=18750 33140 0 0 $X=18670 $Y=32890
X173 35 M2_M1_CDNS_7656633918028 $T=18750 34600 0 0 $X=18670 $Y=34350
X174 35 M2_M1_CDNS_7656633918028 $T=18750 37680 0 0 $X=18670 $Y=37430
X175 35 M2_M1_CDNS_7656633918028 $T=18750 39140 0 0 $X=18670 $Y=38890
X176 35 M2_M1_CDNS_7656633918028 $T=18750 42220 0 0 $X=18670 $Y=41970
X177 35 M2_M1_CDNS_7656633918028 $T=18750 43680 0 0 $X=18670 $Y=43430
X178 35 M2_M1_CDNS_7656633918028 $T=18750 46750 0 0 $X=18670 $Y=46500
X179 35 M2_M1_CDNS_7656633918028 $T=18750 48210 0 0 $X=18670 $Y=47960
X180 44 M2_M1_CDNS_7656633918028 $T=23840 31230 0 0 $X=23760 $Y=30980
X181 44 M2_M1_CDNS_7656633918028 $T=23840 33140 0 0 $X=23760 $Y=32890
X182 44 M2_M1_CDNS_7656633918028 $T=23840 34600 0 0 $X=23760 $Y=34350
X183 44 M2_M1_CDNS_7656633918028 $T=23840 37680 0 0 $X=23760 $Y=37430
X184 44 M2_M1_CDNS_7656633918028 $T=23840 39140 0 0 $X=23760 $Y=38890
X185 44 M2_M1_CDNS_7656633918028 $T=23840 42220 0 0 $X=23760 $Y=41970
X186 44 M2_M1_CDNS_7656633918028 $T=23840 43680 0 0 $X=23760 $Y=43430
X187 44 M2_M1_CDNS_7656633918028 $T=23840 46750 0 0 $X=23760 $Y=46500
X188 44 M2_M1_CDNS_7656633918028 $T=23840 48210 0 0 $X=23760 $Y=47960
X189 53 M2_M1_CDNS_7656633918028 $T=28730 31230 0 0 $X=28650 $Y=30980
X190 53 M2_M1_CDNS_7656633918028 $T=28730 33140 0 0 $X=28650 $Y=32890
X191 53 M2_M1_CDNS_7656633918028 $T=28730 34600 0 0 $X=28650 $Y=34350
X192 53 M2_M1_CDNS_7656633918028 $T=28730 37680 0 0 $X=28650 $Y=37430
X193 53 M2_M1_CDNS_7656633918028 $T=28730 39140 0 0 $X=28650 $Y=38890
X194 53 M2_M1_CDNS_7656633918028 $T=28730 42220 0 0 $X=28650 $Y=41970
X195 53 M2_M1_CDNS_7656633918028 $T=28730 43680 0 0 $X=28650 $Y=43430
X196 53 M2_M1_CDNS_7656633918028 $T=28730 46750 0 0 $X=28650 $Y=46500
X197 53 M2_M1_CDNS_7656633918028 $T=28730 48210 0 0 $X=28650 $Y=47960
X198 62 M2_M1_CDNS_7656633918028 $T=33970 31230 0 0 $X=33890 $Y=30980
X199 62 M2_M1_CDNS_7656633918028 $T=33970 33140 0 0 $X=33890 $Y=32890
X200 62 M2_M1_CDNS_7656633918028 $T=33970 34600 0 0 $X=33890 $Y=34350
X201 62 M2_M1_CDNS_7656633918028 $T=33970 37680 0 0 $X=33890 $Y=37430
X202 62 M2_M1_CDNS_7656633918028 $T=33970 39140 0 0 $X=33890 $Y=38890
X203 62 M2_M1_CDNS_7656633918028 $T=33970 42220 0 0 $X=33890 $Y=41970
X204 62 M2_M1_CDNS_7656633918028 $T=33970 43680 0 0 $X=33890 $Y=43430
X205 62 M2_M1_CDNS_7656633918028 $T=33970 46750 0 0 $X=33890 $Y=46500
X206 62 M2_M1_CDNS_7656633918028 $T=33970 48210 0 0 $X=33890 $Y=47960
X207 71 M2_M1_CDNS_7656633918028 $T=39020 31230 0 0 $X=38940 $Y=30980
X208 71 M2_M1_CDNS_7656633918028 $T=39020 33140 0 0 $X=38940 $Y=32890
X209 71 M2_M1_CDNS_7656633918028 $T=39020 34600 0 0 $X=38940 $Y=34350
X210 71 M2_M1_CDNS_7656633918028 $T=39020 37680 0 0 $X=38940 $Y=37430
X211 71 M2_M1_CDNS_7656633918028 $T=39020 39140 0 0 $X=38940 $Y=38890
X212 71 M2_M1_CDNS_7656633918028 $T=39020 42220 0 0 $X=38940 $Y=41970
X213 71 M2_M1_CDNS_7656633918028 $T=39020 43680 0 0 $X=38940 $Y=43430
X214 71 M2_M1_CDNS_7656633918028 $T=39020 46750 0 0 $X=38940 $Y=46500
X215 71 M2_M1_CDNS_7656633918028 $T=39020 48210 0 0 $X=38940 $Y=47960
X216 1 2 10 11 19 90 154 AND $T=2730 30830 1 0 $X=3800 $Y=31540
X217 1 3 10 11 20 89 153 AND $T=2730 36910 0 0 $X=3800 $Y=33810
X218 1 4 10 11 12 88 152 AND $T=2730 35370 1 0 $X=3800 $Y=36080
X219 1 5 10 11 13 87 151 AND $T=2730 41450 0 0 $X=3800 $Y=38350
X220 1 6 10 11 14 86 150 AND $T=2730 39910 1 0 $X=3800 $Y=40620
X221 1 7 10 11 15 85 149 AND $T=2730 45990 0 0 $X=3800 $Y=42890
X222 1 8 10 11 16 84 148 AND $T=2730 44450 1 0 $X=3800 $Y=45160
X223 1 9 10 11 17 83 147 AND $T=2730 50530 0 0 $X=3800 $Y=47430
X224 18 2 10 11 27 98 162 AND $T=7940 30820 1 0 $X=9010 $Y=31530
X225 18 3 10 11 28 97 161 AND $T=7940 36900 0 0 $X=9010 $Y=33800
X226 18 4 10 11 29 96 160 AND $T=7940 35370 1 0 $X=9010 $Y=36080
X227 18 5 10 11 21 95 159 AND $T=7940 41450 0 0 $X=9010 $Y=38350
X228 18 6 10 11 22 94 158 AND $T=7940 39910 1 0 $X=9010 $Y=40620
X229 18 7 10 11 23 93 157 AND $T=7940 45990 0 0 $X=9010 $Y=42890
X230 18 8 10 11 24 92 156 AND $T=7940 44450 1 0 $X=9010 $Y=45160
X231 18 9 10 11 25 91 155 AND $T=7940 50530 0 0 $X=9010 $Y=47430
X232 26 2 10 11 36 106 170 AND $T=12940 30820 1 0 $X=14010 $Y=31530
X233 26 3 10 11 37 105 169 AND $T=12940 36900 0 0 $X=14010 $Y=33800
X234 26 4 10 11 38 104 168 AND $T=12940 35370 1 0 $X=14010 $Y=36080
X235 26 5 10 11 30 103 167 AND $T=12940 41450 0 0 $X=14010 $Y=38350
X236 26 6 10 11 31 102 166 AND $T=12940 39910 1 0 $X=14010 $Y=40620
X237 26 7 10 11 32 101 165 AND $T=12940 45990 0 0 $X=14010 $Y=42890
X238 26 8 10 11 33 100 164 AND $T=12940 44450 1 0 $X=14010 $Y=45160
X239 26 9 10 11 34 99 163 AND $T=12940 50530 0 0 $X=14010 $Y=47430
X240 35 2 10 11 45 114 178 AND $T=18070 30820 1 0 $X=19140 $Y=31530
X241 35 3 10 11 46 113 177 AND $T=18070 36900 0 0 $X=19140 $Y=33800
X242 35 4 10 11 47 112 176 AND $T=18070 35370 1 0 $X=19140 $Y=36080
X243 35 5 10 11 39 111 175 AND $T=18070 41450 0 0 $X=19140 $Y=38350
X244 35 6 10 11 40 110 174 AND $T=18070 39910 1 0 $X=19140 $Y=40620
X245 35 7 10 11 41 109 173 AND $T=18070 45990 0 0 $X=19140 $Y=42890
X246 35 8 10 11 42 108 172 AND $T=18070 44450 1 0 $X=19140 $Y=45160
X247 35 9 10 11 43 107 171 AND $T=18070 50530 0 0 $X=19140 $Y=47430
X248 44 2 10 11 54 122 186 AND $T=23140 30820 1 0 $X=24210 $Y=31530
X249 44 3 10 11 55 121 185 AND $T=23140 36900 0 0 $X=24210 $Y=33800
X250 44 4 10 11 56 120 184 AND $T=23140 35370 1 0 $X=24210 $Y=36080
X251 44 5 10 11 48 119 183 AND $T=23140 41450 0 0 $X=24210 $Y=38350
X252 44 6 10 11 49 118 182 AND $T=23140 39910 1 0 $X=24210 $Y=40620
X253 44 7 10 11 50 117 181 AND $T=23140 45990 0 0 $X=24210 $Y=42890
X254 44 8 10 11 51 116 180 AND $T=23140 44450 1 0 $X=24210 $Y=45160
X255 44 9 10 11 52 115 179 AND $T=23140 50530 0 0 $X=24210 $Y=47430
X256 53 2 10 11 63 130 194 AND $T=28010 30820 1 0 $X=29080 $Y=31530
X257 53 3 10 11 64 129 193 AND $T=28010 36900 0 0 $X=29080 $Y=33800
X258 53 4 10 11 65 128 192 AND $T=28010 35370 1 0 $X=29080 $Y=36080
X259 53 5 10 11 57 127 191 AND $T=28010 41450 0 0 $X=29080 $Y=38350
X260 53 6 10 11 58 126 190 AND $T=28010 39910 1 0 $X=29080 $Y=40620
X261 53 7 10 11 59 125 189 AND $T=28010 45990 0 0 $X=29080 $Y=42890
X262 53 8 10 11 60 124 188 AND $T=28010 44450 1 0 $X=29080 $Y=45160
X263 53 9 10 11 61 123 187 AND $T=28010 50530 0 0 $X=29080 $Y=47430
X264 62 2 10 11 72 138 202 AND $T=33230 30830 1 0 $X=34300 $Y=31540
X265 62 3 10 11 73 137 201 AND $T=33230 36900 0 0 $X=34300 $Y=33800
X266 62 4 10 11 74 136 200 AND $T=33230 35370 1 0 $X=34300 $Y=36080
X267 62 5 10 11 66 135 199 AND $T=33230 41450 0 0 $X=34300 $Y=38350
X268 62 6 10 11 67 134 198 AND $T=33230 39910 1 0 $X=34300 $Y=40620
X269 62 7 10 11 68 133 197 AND $T=33230 45990 0 0 $X=34300 $Y=42890
X270 62 8 10 11 69 132 196 AND $T=33230 44450 1 0 $X=34300 $Y=45160
X271 62 9 10 11 70 131 195 AND $T=33230 50530 0 0 $X=34300 $Y=47430
X272 71 2 10 11 80 146 210 AND $T=38250 30830 1 0 $X=39320 $Y=31540
X273 71 3 10 11 81 145 209 AND $T=38250 36910 0 0 $X=39320 $Y=33810
X274 71 4 10 11 82 144 208 AND $T=38250 35370 1 0 $X=39320 $Y=36080
X275 71 5 10 11 75 143 207 AND $T=38250 41450 0 0 $X=39320 $Y=38350
X276 71 6 10 11 76 142 206 AND $T=38250 39910 1 0 $X=39320 $Y=40620
X277 71 7 10 11 77 141 205 AND $T=38250 45990 0 0 $X=39320 $Y=42890
X278 71 8 10 11 78 140 204 AND $T=38250 44450 1 0 $X=39320 $Y=45160
X279 71 9 10 11 79 139 203 AND $T=38250 50530 0 0 $X=39320 $Y=47430
X280 17 16 15 14 13 12 20 19 MASCO__Y1 $T=4320 31030 0 0 $X=4320 $Y=31030
X281 25 24 23 22 21 29 28 27 MASCO__Y1 $T=9530 31030 0 0 $X=9530 $Y=31030
X282 34 33 32 31 30 38 37 36 MASCO__Y1 $T=14515 31030 0 0 $X=14515 $Y=31030
X283 43 42 41 40 39 47 46 45 MASCO__Y1 $T=19655 31030 0 0 $X=19655 $Y=31030
X284 52 51 50 49 48 56 55 54 MASCO__Y1 $T=24735 31030 0 0 $X=24735 $Y=31030
X285 61 60 59 58 57 65 64 63 MASCO__Y1 $T=29595 31030 0 0 $X=29595 $Y=31030
X286 70 69 68 67 66 74 73 72 MASCO__Y1 $T=34815 31030 0 0 $X=34815 $Y=31030
X287 79 78 77 76 75 82 81 80 MASCO__Y1 $T=39840 31030 0 0 $X=39840 $Y=31030
X288 17 16 15 14 13 12 20 19 MASCO__Y2 $T=4320 31030 0 0 $X=4320 $Y=31030
X289 25 24 23 22 21 29 28 27 MASCO__Y2 $T=9530 31030 0 0 $X=9530 $Y=31030
X290 34 33 32 31 30 38 37 36 MASCO__Y2 $T=14515 31030 0 0 $X=14515 $Y=31030
X291 43 42 41 40 39 47 46 45 MASCO__Y2 $T=19655 31030 0 0 $X=19655 $Y=31030
X292 52 51 50 49 48 56 55 54 MASCO__Y2 $T=24735 31030 0 0 $X=24735 $Y=31030
X293 61 60 59 58 57 65 64 63 MASCO__Y2 $T=29595 31030 0 0 $X=29595 $Y=31030
X294 70 69 68 67 66 74 73 72 MASCO__Y2 $T=34815 31030 0 0 $X=34815 $Y=31030
X295 79 78 77 76 75 82 81 80 MASCO__Y2 $T=39840 31030 0 0 $X=39840 $Y=31030
M0 154 2 90 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=33350 $dt=0
M1 153 3 89 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=34150 $dt=0
M2 152 4 88 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=37890 $dt=0
M3 151 5 87 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=38690 $dt=0
M4 150 6 86 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=42430 $dt=0
M5 149 7 85 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=43230 $dt=0
M6 148 8 84 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=46970 $dt=0
M7 147 9 83 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4660 $Y=47770 $dt=0
M8 11 1 154 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=33350 $dt=0
M9 11 1 153 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=34150 $dt=0
M10 11 1 152 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=37890 $dt=0
M11 11 1 151 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=38690 $dt=0
M12 11 1 150 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=42430 $dt=0
M13 11 1 149 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=43230 $dt=0
M14 11 1 148 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=46970 $dt=0
M15 11 1 147 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=4870 $Y=47770 $dt=0
M16 19 90 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=33360 $dt=0
M17 20 89 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=34140 $dt=0
M18 12 88 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=37900 $dt=0
M19 13 87 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=38680 $dt=0
M20 14 86 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=42440 $dt=0
M21 15 85 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=43220 $dt=0
M22 16 84 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=46980 $dt=0
M23 17 83 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=7290 $Y=47760 $dt=0
M24 162 2 98 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=33340 $dt=0
M25 161 3 97 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=34140 $dt=0
M26 160 4 96 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=37890 $dt=0
M27 159 5 95 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=38690 $dt=0
M28 158 6 94 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=42430 $dt=0
M29 157 7 93 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=43230 $dt=0
M30 156 8 92 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=46970 $dt=0
M31 155 9 91 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=9870 $Y=47770 $dt=0
M32 11 18 162 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=33340 $dt=0
M33 11 18 161 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=34140 $dt=0
M34 11 18 160 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=37890 $dt=0
M35 11 18 159 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=38690 $dt=0
M36 11 18 158 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=42430 $dt=0
M37 11 18 157 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=43230 $dt=0
M38 11 18 156 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=46970 $dt=0
M39 11 18 155 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=10080 $Y=47770 $dt=0
M40 27 98 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=33350 $dt=0
M41 28 97 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=34130 $dt=0
M42 29 96 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=37900 $dt=0
M43 21 95 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=38680 $dt=0
M44 22 94 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=42440 $dt=0
M45 23 93 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=43220 $dt=0
M46 24 92 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=46980 $dt=0
M47 25 91 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=12500 $Y=47760 $dt=0
M48 170 2 106 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=33340 $dt=0
M49 169 3 105 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=34140 $dt=0
M50 168 4 104 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=37890 $dt=0
M51 167 5 103 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=38690 $dt=0
M52 166 6 102 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=42430 $dt=0
M53 165 7 101 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=43230 $dt=0
M54 164 8 100 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=46970 $dt=0
M55 163 9 99 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=14870 $Y=47770 $dt=0
M56 11 26 170 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=33340 $dt=0
M57 11 26 169 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=34140 $dt=0
M58 11 26 168 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=37890 $dt=0
M59 11 26 167 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=38690 $dt=0
M60 11 26 166 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=42430 $dt=0
M61 11 26 165 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=43230 $dt=0
M62 11 26 164 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=46970 $dt=0
M63 11 26 163 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=15080 $Y=47770 $dt=0
M64 36 106 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=33350 $dt=0
M65 37 105 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=34130 $dt=0
M66 38 104 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=37900 $dt=0
M67 30 103 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=38680 $dt=0
M68 31 102 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=42440 $dt=0
M69 32 101 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=43220 $dt=0
M70 33 100 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=46980 $dt=0
M71 34 99 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=17500 $Y=47760 $dt=0
M72 178 2 114 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=33340 $dt=0
M73 177 3 113 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=34140 $dt=0
M74 176 4 112 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=37890 $dt=0
M75 175 5 111 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=38690 $dt=0
M76 174 6 110 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=42430 $dt=0
M77 173 7 109 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=43230 $dt=0
M78 172 8 108 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=46970 $dt=0
M79 171 9 107 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20000 $Y=47770 $dt=0
M80 11 35 178 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=33340 $dt=0
M81 11 35 177 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=34140 $dt=0
M82 11 35 176 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=37890 $dt=0
M83 11 35 175 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=38690 $dt=0
M84 11 35 174 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=42430 $dt=0
M85 11 35 173 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=43230 $dt=0
M86 11 35 172 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=46970 $dt=0
M87 11 35 171 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=20210 $Y=47770 $dt=0
M88 45 114 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=33350 $dt=0
M89 46 113 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=34130 $dt=0
M90 47 112 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=37900 $dt=0
M91 39 111 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=38680 $dt=0
M92 40 110 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=42440 $dt=0
M93 41 109 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=43220 $dt=0
M94 42 108 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=46980 $dt=0
M95 43 107 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=22630 $Y=47760 $dt=0
M96 186 2 122 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=33340 $dt=0
M97 185 3 121 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=34140 $dt=0
M98 184 4 120 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=37890 $dt=0
M99 183 5 119 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=38690 $dt=0
M100 182 6 118 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=42430 $dt=0
M101 181 7 117 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=43230 $dt=0
M102 180 8 116 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=46970 $dt=0
M103 179 9 115 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25070 $Y=47770 $dt=0
M104 11 44 186 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=33340 $dt=0
M105 11 44 185 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=34140 $dt=0
M106 11 44 184 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=37890 $dt=0
M107 11 44 183 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=38690 $dt=0
M108 11 44 182 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=42430 $dt=0
M109 11 44 181 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=43230 $dt=0
M110 11 44 180 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=46970 $dt=0
M111 11 44 179 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=25280 $Y=47770 $dt=0
M112 54 122 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=33350 $dt=0
M113 55 121 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=34130 $dt=0
M114 56 120 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=37900 $dt=0
M115 48 119 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=38680 $dt=0
M116 49 118 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=42440 $dt=0
M117 50 117 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=43220 $dt=0
M118 51 116 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=46980 $dt=0
M119 52 115 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=27700 $Y=47760 $dt=0
M120 194 2 130 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=33340 $dt=0
M121 193 3 129 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=34140 $dt=0
M122 192 4 128 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=37890 $dt=0
M123 191 5 127 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=38690 $dt=0
M124 190 6 126 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=42430 $dt=0
M125 189 7 125 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=43230 $dt=0
M126 188 8 124 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=46970 $dt=0
M127 187 9 123 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=29940 $Y=47770 $dt=0
M128 11 53 194 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=33340 $dt=0
M129 11 53 193 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=34140 $dt=0
M130 11 53 192 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=37890 $dt=0
M131 11 53 191 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=38690 $dt=0
M132 11 53 190 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=42430 $dt=0
M133 11 53 189 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=43230 $dt=0
M134 11 53 188 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=46970 $dt=0
M135 11 53 187 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=30150 $Y=47770 $dt=0
M136 63 130 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=33350 $dt=0
M137 64 129 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=34130 $dt=0
M138 65 128 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=37900 $dt=0
M139 57 127 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=38680 $dt=0
M140 58 126 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=42440 $dt=0
M141 59 125 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=43220 $dt=0
M142 60 124 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=46980 $dt=0
M143 61 123 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=32570 $Y=47760 $dt=0
M144 202 2 138 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=33350 $dt=0
M145 201 3 137 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35160 $Y=34140 $dt=0
M146 200 4 136 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=37890 $dt=0
M147 199 5 135 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=38690 $dt=0
M148 198 6 134 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=42430 $dt=0
M149 197 7 133 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=43230 $dt=0
M150 196 8 132 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=46970 $dt=0
M151 195 9 131 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35160 $Y=47770 $dt=0
M152 11 62 202 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=33350 $dt=0
M153 11 62 201 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.13128 scb=0.00354568 scc=2.49792e-05 $X=35370 $Y=34140 $dt=0
M154 11 62 200 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=37890 $dt=0
M155 11 62 199 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=38690 $dt=0
M156 11 62 198 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=42430 $dt=0
M157 11 62 197 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=43230 $dt=0
M158 11 62 196 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=46970 $dt=0
M159 11 62 195 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=35370 $Y=47770 $dt=0
M160 72 138 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=33360 $dt=0
M161 73 137 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.06655 scb=0.00341969 scc=2.28395e-05 $X=37790 $Y=34130 $dt=0
M162 74 136 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=37900 $dt=0
M163 66 135 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=38680 $dt=0
M164 67 134 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=42440 $dt=0
M165 68 133 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=43220 $dt=0
M166 69 132 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=46980 $dt=0
M167 70 131 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=37790 $Y=47760 $dt=0
M168 210 2 146 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=33350 $dt=0
M169 209 3 145 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=34150 $dt=0
M170 208 4 144 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=37890 $dt=0
M171 207 5 143 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=38690 $dt=0
M172 206 6 142 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=42430 $dt=0
M173 205 7 141 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=43230 $dt=0
M174 204 8 140 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=46970 $dt=0
M175 203 9 139 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40180 $Y=47770 $dt=0
M176 11 71 210 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=33350 $dt=0
M177 11 71 209 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=34150 $dt=0
M178 11 71 208 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=37890 $dt=0
M179 11 71 207 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=38690 $dt=0
M180 11 71 206 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=42430 $dt=0
M181 11 71 205 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=43230 $dt=0
M182 11 71 204 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=46970 $dt=0
M183 11 71 203 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.11756 scb=0.00354063 scc=2.49777e-05 $X=40390 $Y=47770 $dt=0
M184 80 146 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=33360 $dt=0
M185 81 145 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=34140 $dt=0
M186 82 144 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=37900 $dt=0
M187 75 143 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=38680 $dt=0
M188 76 142 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=42440 $dt=0
M189 77 141 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=43220 $dt=0
M190 78 140 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=46980 $dt=0
M191 79 139 11 11 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=7.05259 scb=0.00341442 scc=2.28378e-05 $X=42810 $Y=47760 $dt=0
M192 90 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=31910 $dt=1
M193 89 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=35590 $dt=1
M194 88 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=36450 $dt=1
M195 87 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40130 $dt=1
M196 86 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=40990 $dt=1
M197 85 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=44670 $dt=1
M198 84 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=4660 $Y=45530 $dt=1
M199 83 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=4660 $Y=49210 $dt=1
M200 10 1 90 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=31910 $dt=1
M201 10 1 89 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=35590 $dt=1
M202 10 1 88 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=36450 $dt=1
M203 10 1 87 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40130 $dt=1
M204 10 1 86 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=40990 $dt=1
M205 10 1 85 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=44670 $dt=1
M206 10 1 84 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=5070 $Y=45530 $dt=1
M207 10 1 83 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=5070 $Y=49210 $dt=1
M208 19 90 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=31860 $dt=1
M209 20 89 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=35400 $dt=1
M210 12 88 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=36400 $dt=1
M211 13 87 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=39940 $dt=1
M212 14 86 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=40940 $dt=1
M213 15 85 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=44480 $dt=1
M214 16 84 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=7290 $Y=45480 $dt=1
M215 17 83 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=7290 $Y=49020 $dt=1
M216 98 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=31900 $dt=1
M217 97 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=35580 $dt=1
M218 96 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=9870 $Y=36450 $dt=1
M219 95 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40130 $dt=1
M220 94 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=40990 $dt=1
M221 93 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=44670 $dt=1
M222 92 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=9870 $Y=45530 $dt=1
M223 91 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=9870 $Y=49210 $dt=1
M224 10 18 98 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=31900 $dt=1
M225 10 18 97 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=35580 $dt=1
M226 10 18 96 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=10280 $Y=36450 $dt=1
M227 10 18 95 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40130 $dt=1
M228 10 18 94 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=40990 $dt=1
M229 10 18 93 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=44670 $dt=1
M230 10 18 92 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=10280 $Y=45530 $dt=1
M231 10 18 91 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=10280 $Y=49210 $dt=1
M232 27 98 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=31850 $dt=1
M233 28 97 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=35390 $dt=1
M234 29 96 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=12500 $Y=36400 $dt=1
M235 21 95 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=39940 $dt=1
M236 22 94 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=40940 $dt=1
M237 23 93 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=44480 $dt=1
M238 24 92 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=12500 $Y=45480 $dt=1
M239 25 91 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=12500 $Y=49020 $dt=1
M240 106 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=31900 $dt=1
M241 105 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=35580 $dt=1
M242 104 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=14870 $Y=36450 $dt=1
M243 103 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40130 $dt=1
M244 102 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=40990 $dt=1
M245 101 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=44670 $dt=1
M246 100 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=14870 $Y=45530 $dt=1
M247 99 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14870 $Y=49210 $dt=1
M248 10 26 106 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=31900 $dt=1
M249 10 26 105 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=35580 $dt=1
M250 10 26 104 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=15280 $Y=36450 $dt=1
M251 10 26 103 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40130 $dt=1
M252 10 26 102 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=40990 $dt=1
M253 10 26 101 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=44670 $dt=1
M254 10 26 100 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=15280 $Y=45530 $dt=1
M255 10 26 99 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=15280 $Y=49210 $dt=1
M256 36 106 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=31850 $dt=1
M257 37 105 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=35390 $dt=1
M258 38 104 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=17500 $Y=36400 $dt=1
M259 30 103 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=39940 $dt=1
M260 31 102 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=40940 $dt=1
M261 32 101 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=44480 $dt=1
M262 33 100 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=17500 $Y=45480 $dt=1
M263 34 99 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17500 $Y=49020 $dt=1
M264 114 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=31900 $dt=1
M265 113 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=35580 $dt=1
M266 112 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=20000 $Y=36450 $dt=1
M267 111 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40130 $dt=1
M268 110 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=40990 $dt=1
M269 109 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=44670 $dt=1
M270 108 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=20000 $Y=45530 $dt=1
M271 107 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=20000 $Y=49210 $dt=1
M272 10 35 114 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=31900 $dt=1
M273 10 35 113 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=35580 $dt=1
M274 10 35 112 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=20410 $Y=36450 $dt=1
M275 10 35 111 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40130 $dt=1
M276 10 35 110 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=40990 $dt=1
M277 10 35 109 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=44670 $dt=1
M278 10 35 108 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=20410 $Y=45530 $dt=1
M279 10 35 107 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20410 $Y=49210 $dt=1
M280 45 114 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=31850 $dt=1
M281 46 113 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=35390 $dt=1
M282 47 112 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=22630 $Y=36400 $dt=1
M283 39 111 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=39940 $dt=1
M284 40 110 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=40940 $dt=1
M285 41 109 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=44480 $dt=1
M286 42 108 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=22630 $Y=45480 $dt=1
M287 43 107 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22630 $Y=49020 $dt=1
M288 122 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=31900 $dt=1
M289 121 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=35580 $dt=1
M290 120 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=25070 $Y=36450 $dt=1
M291 119 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40130 $dt=1
M292 118 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=40990 $dt=1
M293 117 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=44670 $dt=1
M294 116 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=25070 $Y=45530 $dt=1
M295 115 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=25070 $Y=49210 $dt=1
M296 10 44 122 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=31900 $dt=1
M297 10 44 121 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=35580 $dt=1
M298 10 44 120 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=25480 $Y=36450 $dt=1
M299 10 44 119 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40130 $dt=1
M300 10 44 118 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=40990 $dt=1
M301 10 44 117 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=44670 $dt=1
M302 10 44 116 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=25480 $Y=45530 $dt=1
M303 10 44 115 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=25480 $Y=49210 $dt=1
M304 54 122 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=31850 $dt=1
M305 55 121 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=35390 $dt=1
M306 56 120 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=27700 $Y=36400 $dt=1
M307 48 119 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=39940 $dt=1
M308 49 118 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=40940 $dt=1
M309 50 117 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=44480 $dt=1
M310 51 116 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=27700 $Y=45480 $dt=1
M311 52 115 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27700 $Y=49020 $dt=1
M312 130 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=31900 $dt=1
M313 129 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=35580 $dt=1
M314 128 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=29940 $Y=36450 $dt=1
M315 127 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40130 $dt=1
M316 126 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=40990 $dt=1
M317 125 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=44670 $dt=1
M318 124 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=29940 $Y=45530 $dt=1
M319 123 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=29940 $Y=49210 $dt=1
M320 10 53 130 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=31900 $dt=1
M321 10 53 129 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=35580 $dt=1
M322 10 53 128 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=30350 $Y=36450 $dt=1
M323 10 53 127 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40130 $dt=1
M324 10 53 126 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=40990 $dt=1
M325 10 53 125 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=44670 $dt=1
M326 10 53 124 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=30350 $Y=45530 $dt=1
M327 10 53 123 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=30350 $Y=49210 $dt=1
M328 63 130 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=31850 $dt=1
M329 64 129 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=35390 $dt=1
M330 65 128 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=32570 $Y=36400 $dt=1
M331 57 127 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=39940 $dt=1
M332 58 126 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=40940 $dt=1
M333 59 125 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=44480 $dt=1
M334 60 124 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=32570 $Y=45480 $dt=1
M335 61 123 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=32570 $Y=49020 $dt=1
M336 138 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=31910 $dt=1
M337 137 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=35580 $dt=1
M338 136 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.444 scb=0.0358776 scc=0.00356009 $X=35160 $Y=36450 $dt=1
M339 135 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40130 $dt=1
M340 134 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=40990 $dt=1
M341 133 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=44670 $dt=1
M342 132 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=35160 $Y=45530 $dt=1
M343 131 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=35160 $Y=49210 $dt=1
M344 10 62 138 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=31910 $dt=1
M345 10 62 137 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=35580 $dt=1
M346 10 62 136 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.9145 scb=0.0281383 scc=0.00330319 $X=35570 $Y=36450 $dt=1
M347 10 62 135 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40130 $dt=1
M348 10 62 134 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=40990 $dt=1
M349 10 62 133 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=44670 $dt=1
M350 10 62 132 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=35570 $Y=45530 $dt=1
M351 10 62 131 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=35570 $Y=49210 $dt=1
M352 72 138 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=31860 $dt=1
M353 73 137 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=35390 $dt=1
M354 74 136 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1193 scb=0.0532463 scc=0.00937005 $X=37790 $Y=36400 $dt=1
M355 66 135 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=39940 $dt=1
M356 67 134 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=40940 $dt=1
M357 68 133 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=44480 $dt=1
M358 69 132 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=37790 $Y=45480 $dt=1
M359 70 131 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=37790 $Y=49020 $dt=1
M360 146 2 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=31910 $dt=1
M361 145 3 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=35590 $dt=1
M362 144 4 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=36450 $dt=1
M363 143 5 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40130 $dt=1
M364 142 6 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=40990 $dt=1
M365 141 7 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=44670 $dt=1
M366 140 8 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=34.4815 scb=0.0359214 scc=0.00356026 $X=40180 $Y=45530 $dt=1
M367 139 9 10 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=40180 $Y=49210 $dt=1
M368 10 71 146 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=31910 $dt=1
M369 10 71 145 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=35590 $dt=1
M370 10 71 144 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=36450 $dt=1
M371 10 71 143 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40130 $dt=1
M372 10 71 142 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=40990 $dt=1
M373 10 71 141 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=44670 $dt=1
M374 10 71 140 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=29.952 scb=0.0281822 scc=0.00330336 $X=40590 $Y=45530 $dt=1
M375 10 71 139 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=40590 $Y=49210 $dt=1
M376 80 146 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=31860 $dt=1
M377 81 145 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=35400 $dt=1
M378 82 144 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=36400 $dt=1
M379 75 143 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=39940 $dt=1
M380 76 142 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=40940 $dt=1
M381 77 141 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=44480 $dt=1
M382 78 140 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=79.1528 scb=0.0532831 scc=0.0093702 $X=42810 $Y=45480 $dt=1
M383 79 139 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=42810 $Y=49020 $dt=1
.ends WallaceMultiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: Diver                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt Diver 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
X0 1 M1_PO_CDNS_7656633918062 $T=1260 -2440 0 0 $X=1160 $Y=-2560
X1 5 M1_PO_CDNS_7656633918062 $T=2200 -2440 0 0 $X=2100 $Y=-2560
X2 2 2 1 5 3 pmos1v_CDNS_765663391806 $T=1340 -2060 0 0 $X=920 $Y=-2260
X3 2 2 5 4 3 pmos1v_CDNS_765663391806 $T=2270 -2060 0 0 $X=1850 $Y=-2260
X4 3 3 1 5 nmos1v_CDNS_765663391807 $T=1340 -3070 0 0 $X=920 $Y=-3630
X5 3 3 5 4 nmos1v_CDNS_765663391807 $T=2270 -3070 0 0 $X=1850 $Y=-3630
.ends Diver

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MAC                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MAC 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96
** N=288 EP=96 FDC=570
X0 52 M4_M3_CDNS_765663391804 $T=57860 9670 0 90 $X=57730 $Y=9590
X1 5 M2_M1_CDNS_765663391809 $T=9840 3330 0 0 $X=9760 $Y=3080
X2 53 M4_M3_CDNS_7656633918010 $T=150 23850 0 0 $X=70 $Y=23600
X3 54 M4_M3_CDNS_7656633918010 $T=5940 23850 0 0 $X=5860 $Y=23600
X4 55 M4_M3_CDNS_7656633918010 $T=16170 2650 0 0 $X=16090 $Y=2400
X5 56 M4_M3_CDNS_7656633918010 $T=16170 23850 0 0 $X=16090 $Y=23600
X6 57 M4_M3_CDNS_7656633918010 $T=21750 2650 0 0 $X=21670 $Y=2400
X7 58 M4_M3_CDNS_7656633918010 $T=21750 23850 0 0 $X=21670 $Y=23600
X8 59 M4_M3_CDNS_7656633918010 $T=26890 2650 0 0 $X=26810 $Y=2400
X9 60 M4_M3_CDNS_7656633918010 $T=26890 23850 0 0 $X=26810 $Y=23600
X10 61 M4_M3_CDNS_7656633918010 $T=32670 2650 0 0 $X=32590 $Y=2400
X11 62 M4_M3_CDNS_7656633918010 $T=32670 23850 0 0 $X=32590 $Y=23600
X12 63 M4_M3_CDNS_7656633918010 $T=40090 2650 0 0 $X=40010 $Y=2400
X13 33 M4_M3_CDNS_7656633918010 $T=40090 23850 0 0 $X=40010 $Y=23600
X14 64 M4_M3_CDNS_7656633918010 $T=48440 2650 0 0 $X=48360 $Y=2400
X15 33 M4_M3_CDNS_7656633918010 $T=48440 23850 0 0 $X=48360 $Y=23600
X16 33 M4_M3_CDNS_7656633918010 $T=53580 23850 0 0 $X=53500 $Y=23600
X17 53 M3_M2_CDNS_7656633918011 $T=150 23850 0 0 $X=70 $Y=23600
X18 54 M3_M2_CDNS_7656633918011 $T=5940 23850 0 0 $X=5860 $Y=23600
X19 5 M3_M2_CDNS_7656633918011 $T=9840 3330 0 0 $X=9760 $Y=3080
X20 55 M3_M2_CDNS_7656633918011 $T=16170 2650 0 0 $X=16090 $Y=2400
X21 56 M3_M2_CDNS_7656633918011 $T=16170 23850 0 0 $X=16090 $Y=23600
X22 57 M3_M2_CDNS_7656633918011 $T=21750 2650 0 0 $X=21670 $Y=2400
X23 58 M3_M2_CDNS_7656633918011 $T=21750 23850 0 0 $X=21670 $Y=23600
X24 59 M3_M2_CDNS_7656633918011 $T=26890 2650 0 0 $X=26810 $Y=2400
X25 60 M3_M2_CDNS_7656633918011 $T=26890 23850 0 0 $X=26810 $Y=23600
X26 61 M3_M2_CDNS_7656633918011 $T=32670 2650 0 0 $X=32590 $Y=2400
X27 62 M3_M2_CDNS_7656633918011 $T=32670 23850 0 0 $X=32590 $Y=23600
X28 63 M3_M2_CDNS_7656633918011 $T=40090 2650 0 0 $X=40010 $Y=2400
X29 33 M3_M2_CDNS_7656633918011 $T=40090 23850 0 0 $X=40010 $Y=23600
X30 64 M3_M2_CDNS_7656633918011 $T=48440 2650 0 0 $X=48360 $Y=2400
X31 33 M3_M2_CDNS_7656633918011 $T=48440 23850 0 0 $X=48360 $Y=23600
X32 33 M3_M2_CDNS_7656633918011 $T=53580 23850 0 0 $X=53500 $Y=23600
X33 1 M2_M1_CDNS_7656633918020 $T=4820 41440 0 0 $X=4740 $Y=41310
X34 8 M2_M1_CDNS_7656633918020 $T=13610 20240 0 0 $X=13530 $Y=20110
X35 9 M2_M1_CDNS_7656633918020 $T=13610 41440 0 0 $X=13530 $Y=41310
X36 14 M2_M1_CDNS_7656633918020 $T=19200 20240 0 0 $X=19120 $Y=20110
X37 15 M2_M1_CDNS_7656633918020 $T=19200 41440 0 0 $X=19120 $Y=41310
X38 22 M2_M1_CDNS_7656633918020 $T=31060 20240 0 0 $X=30980 $Y=20110
X39 23 M2_M1_CDNS_7656633918020 $T=31060 41440 0 0 $X=30980 $Y=41310
X40 24 M2_M1_CDNS_7656633918020 $T=31510 20240 0 0 $X=31430 $Y=20110
X41 25 M2_M1_CDNS_7656633918020 $T=31510 41440 0 0 $X=31430 $Y=41310
X42 32 M2_M1_CDNS_7656633918020 $T=40300 20240 0 0 $X=40220 $Y=20110
X43 33 M2_M1_CDNS_7656633918020 $T=40300 41440 0 0 $X=40220 $Y=41310
X44 38 M2_M1_CDNS_7656633918020 $T=45890 20240 0 0 $X=45810 $Y=20110
X45 39 M2_M1_CDNS_7656633918020 $T=45890 41440 0 0 $X=45810 $Y=41310
X46 48 M2_M1_CDNS_7656633918020 $T=57710 20240 0 0 $X=57630 $Y=20110
X47 49 M2_M1_CDNS_7656633918020 $T=57710 41440 0 0 $X=57630 $Y=41310
X48 52 M3_M2_CDNS_7656633918035 $T=560 24410 0 0 $X=480 $Y=24160
X49 65 M3_M2_CDNS_7656633918035 $T=9840 24410 0 0 $X=9760 $Y=24160
X50 66 M3_M2_CDNS_7656633918035 $T=17280 3210 0 0 $X=17200 $Y=2960
X51 67 M3_M2_CDNS_7656633918035 $T=17280 24410 0 0 $X=17200 $Y=24160
X52 68 M3_M2_CDNS_7656633918035 $T=22860 3210 0 0 $X=22780 $Y=2960
X53 69 M3_M2_CDNS_7656633918035 $T=22860 24410 0 0 $X=22780 $Y=24160
X54 70 M3_M2_CDNS_7656633918035 $T=27230 3210 0 0 $X=27150 $Y=2960
X55 71 M3_M2_CDNS_7656633918035 $T=27230 24410 0 0 $X=27150 $Y=24160
X56 72 M3_M2_CDNS_7656633918035 $T=36530 3210 0 0 $X=36450 $Y=2960
X57 73 M3_M2_CDNS_7656633918035 $T=36530 24410 0 0 $X=36450 $Y=24160
X58 74 M3_M2_CDNS_7656633918035 $T=43970 3210 0 0 $X=43890 $Y=2960
X59 75 M3_M2_CDNS_7656633918035 $T=43970 24410 0 0 $X=43890 $Y=24160
X60 76 M3_M2_CDNS_7656633918035 $T=49550 3210 0 0 $X=49470 $Y=2960
X61 77 M3_M2_CDNS_7656633918035 $T=49550 24410 0 0 $X=49470 $Y=24160
X62 52 M4_M3_CDNS_7656633918036 $T=560 24410 0 0 $X=480 $Y=24160
X63 5 M4_M3_CDNS_7656633918036 $T=9840 3330 0 0 $X=9760 $Y=3080
X64 65 M4_M3_CDNS_7656633918036 $T=9840 24410 0 0 $X=9760 $Y=24160
X65 66 M4_M3_CDNS_7656633918036 $T=17280 3210 0 0 $X=17200 $Y=2960
X66 67 M4_M3_CDNS_7656633918036 $T=17280 24410 0 0 $X=17200 $Y=24160
X67 68 M4_M3_CDNS_7656633918036 $T=22860 3210 0 0 $X=22780 $Y=2960
X68 69 M4_M3_CDNS_7656633918036 $T=22860 24410 0 0 $X=22780 $Y=24160
X69 70 M4_M3_CDNS_7656633918036 $T=27230 3210 0 0 $X=27150 $Y=2960
X70 71 M4_M3_CDNS_7656633918036 $T=27230 24410 0 0 $X=27150 $Y=24160
X71 72 M4_M3_CDNS_7656633918036 $T=36530 3210 0 0 $X=36450 $Y=2960
X72 73 M4_M3_CDNS_7656633918036 $T=36530 24410 0 0 $X=36450 $Y=24160
X73 74 M4_M3_CDNS_7656633918036 $T=43970 3210 0 0 $X=43890 $Y=2960
X74 75 M4_M3_CDNS_7656633918036 $T=43970 24410 0 0 $X=43890 $Y=24160
X75 76 M4_M3_CDNS_7656633918036 $T=49550 3210 0 0 $X=49470 $Y=2960
X76 77 M4_M3_CDNS_7656633918036 $T=49550 24410 0 0 $X=49470 $Y=24160
X77 53 M5_M4_CDNS_7656633918045 $T=150 23850 0 0 $X=70 $Y=23600
X78 54 M5_M4_CDNS_7656633918045 $T=5940 23850 0 0 $X=5860 $Y=23600
X79 55 M5_M4_CDNS_7656633918045 $T=16170 2650 0 0 $X=16090 $Y=2400
X80 56 M5_M4_CDNS_7656633918045 $T=16170 23850 0 0 $X=16090 $Y=23600
X81 57 M5_M4_CDNS_7656633918045 $T=21750 2650 0 0 $X=21670 $Y=2400
X82 58 M5_M4_CDNS_7656633918045 $T=21750 23850 0 0 $X=21670 $Y=23600
X83 59 M5_M4_CDNS_7656633918045 $T=26890 2650 0 0 $X=26810 $Y=2400
X84 60 M5_M4_CDNS_7656633918045 $T=26890 23850 0 0 $X=26810 $Y=23600
X85 61 M5_M4_CDNS_7656633918045 $T=32670 2650 0 0 $X=32590 $Y=2400
X86 62 M5_M4_CDNS_7656633918045 $T=32670 23850 0 0 $X=32590 $Y=23600
X87 63 M5_M4_CDNS_7656633918045 $T=40090 2650 0 0 $X=40010 $Y=2400
X88 33 M5_M4_CDNS_7656633918045 $T=40090 23850 0 0 $X=40010 $Y=23600
X89 64 M5_M4_CDNS_7656633918045 $T=48440 2650 0 0 $X=48360 $Y=2400
X90 33 M5_M4_CDNS_7656633918045 $T=48440 23850 0 0 $X=48360 $Y=23600
X91 33 M5_M4_CDNS_7656633918045 $T=53580 23850 0 0 $X=53500 $Y=23600
X92 53 M6_M5_CDNS_7656633918053 $T=150 23850 0 0 $X=70 $Y=23600
X93 54 M6_M5_CDNS_7656633918053 $T=5940 23850 0 0 $X=5860 $Y=23600
X94 55 M6_M5_CDNS_7656633918053 $T=16170 2650 0 0 $X=16090 $Y=2400
X95 56 M6_M5_CDNS_7656633918053 $T=16170 23850 0 0 $X=16090 $Y=23600
X96 57 M6_M5_CDNS_7656633918053 $T=21750 2650 0 0 $X=21670 $Y=2400
X97 58 M6_M5_CDNS_7656633918053 $T=21750 23850 0 0 $X=21670 $Y=23600
X98 59 M6_M5_CDNS_7656633918053 $T=26890 2650 0 0 $X=26810 $Y=2400
X99 60 M6_M5_CDNS_7656633918053 $T=26890 23850 0 0 $X=26810 $Y=23600
X100 61 M6_M5_CDNS_7656633918053 $T=32670 2650 0 0 $X=32590 $Y=2400
X101 62 M6_M5_CDNS_7656633918053 $T=32670 23850 0 0 $X=32590 $Y=23600
X102 63 M6_M5_CDNS_7656633918053 $T=40090 2650 0 0 $X=40010 $Y=2400
X103 33 M6_M5_CDNS_7656633918053 $T=40090 23850 0 0 $X=40010 $Y=23600
X104 64 M6_M5_CDNS_7656633918053 $T=48440 2650 0 0 $X=48360 $Y=2400
X105 33 M6_M5_CDNS_7656633918053 $T=48440 23850 0 0 $X=48360 $Y=23600
X106 33 M6_M5_CDNS_7656633918053 $T=53580 23850 0 0 $X=53500 $Y=23600
X107 78 M5_M4_CDNS_7656633918057 $T=9340 41110 0 0 $X=9120 $Y=40860
X108 79 M5_M4_CDNS_7656633918057 $T=18130 19910 0 0 $X=17910 $Y=19660
X109 80 M5_M4_CDNS_7656633918057 $T=18130 41110 0 0 $X=17910 $Y=40860
X110 81 M5_M4_CDNS_7656633918057 $T=23720 19910 0 0 $X=23500 $Y=19660
X111 82 M5_M4_CDNS_7656633918057 $T=23720 41110 0 0 $X=23500 $Y=40860
X112 83 M5_M4_CDNS_7656633918057 $T=26500 19910 0 0 $X=26280 $Y=19660
X113 84 M5_M4_CDNS_7656633918057 $T=26500 41110 0 0 $X=26280 $Y=40860
X114 85 M5_M4_CDNS_7656633918057 $T=36030 19910 0 0 $X=35810 $Y=19660
X115 86 M5_M4_CDNS_7656633918057 $T=36030 41110 0 0 $X=35810 $Y=40860
X116 87 M5_M4_CDNS_7656633918057 $T=44820 19910 0 0 $X=44600 $Y=19660
X117 88 M5_M4_CDNS_7656633918057 $T=44820 41110 0 0 $X=44600 $Y=40860
X118 89 M5_M4_CDNS_7656633918057 $T=50410 19910 0 0 $X=50190 $Y=19660
X119 90 M5_M4_CDNS_7656633918057 $T=50410 41110 0 0 $X=50190 $Y=40860
X120 91 M5_M4_CDNS_7656633918057 $T=53190 19910 0 0 $X=52970 $Y=19660
X121 92 M5_M4_CDNS_7656633918057 $T=53190 41110 0 0 $X=52970 $Y=40860
X122 78 M4_M3_CDNS_7656633918058 $T=9340 41110 0 0 $X=9120 $Y=40860
X123 79 M4_M3_CDNS_7656633918058 $T=18130 19910 0 0 $X=17910 $Y=19660
X124 80 M4_M3_CDNS_7656633918058 $T=18130 41110 0 0 $X=17910 $Y=40860
X125 81 M4_M3_CDNS_7656633918058 $T=23720 19910 0 0 $X=23500 $Y=19660
X126 82 M4_M3_CDNS_7656633918058 $T=23720 41110 0 0 $X=23500 $Y=40860
X127 83 M4_M3_CDNS_7656633918058 $T=26500 19910 0 0 $X=26280 $Y=19660
X128 84 M4_M3_CDNS_7656633918058 $T=26500 41110 0 0 $X=26280 $Y=40860
X129 85 M4_M3_CDNS_7656633918058 $T=36030 19910 0 0 $X=35810 $Y=19660
X130 86 M4_M3_CDNS_7656633918058 $T=36030 41110 0 0 $X=35810 $Y=40860
X131 87 M4_M3_CDNS_7656633918058 $T=44820 19910 0 0 $X=44600 $Y=19660
X132 88 M4_M3_CDNS_7656633918058 $T=44820 41110 0 0 $X=44600 $Y=40860
X133 89 M4_M3_CDNS_7656633918058 $T=50410 19910 0 0 $X=50190 $Y=19660
X134 90 M4_M3_CDNS_7656633918058 $T=50410 41110 0 0 $X=50190 $Y=40860
X135 91 M4_M3_CDNS_7656633918058 $T=53190 19910 0 0 $X=52970 $Y=19660
X136 92 M4_M3_CDNS_7656633918058 $T=53190 41110 0 0 $X=52970 $Y=40860
X137 78 M3_M2_CDNS_7656633918059 $T=9340 41110 0 0 $X=9120 $Y=40860
X138 79 M3_M2_CDNS_7656633918059 $T=18130 19910 0 0 $X=17910 $Y=19660
X139 80 M3_M2_CDNS_7656633918059 $T=18130 41110 0 0 $X=17910 $Y=40860
X140 81 M3_M2_CDNS_7656633918059 $T=23720 19910 0 0 $X=23500 $Y=19660
X141 82 M3_M2_CDNS_7656633918059 $T=23720 41110 0 0 $X=23500 $Y=40860
X142 83 M3_M2_CDNS_7656633918059 $T=26500 19910 0 0 $X=26280 $Y=19660
X143 84 M3_M2_CDNS_7656633918059 $T=26500 41110 0 0 $X=26280 $Y=40860
X144 85 M3_M2_CDNS_7656633918059 $T=36030 19910 0 0 $X=35810 $Y=19660
X145 86 M3_M2_CDNS_7656633918059 $T=36030 41110 0 0 $X=35810 $Y=40860
X146 87 M3_M2_CDNS_7656633918059 $T=44820 19910 0 0 $X=44600 $Y=19660
X147 88 M3_M2_CDNS_7656633918059 $T=44820 41110 0 0 $X=44600 $Y=40860
X148 89 M3_M2_CDNS_7656633918059 $T=50410 19910 0 0 $X=50190 $Y=19660
X149 90 M3_M2_CDNS_7656633918059 $T=50410 41110 0 0 $X=50190 $Y=40860
X150 91 M3_M2_CDNS_7656633918059 $T=53190 19910 0 0 $X=52970 $Y=19660
X151 92 M3_M2_CDNS_7656633918059 $T=53190 41110 0 0 $X=52970 $Y=40860
X152 78 M2_M1_CDNS_7656633918060 $T=9340 41110 0 0 $X=9120 $Y=40860
X153 79 M2_M1_CDNS_7656633918060 $T=18130 19910 0 0 $X=17910 $Y=19660
X154 80 M2_M1_CDNS_7656633918060 $T=18130 41110 0 0 $X=17910 $Y=40860
X155 81 M2_M1_CDNS_7656633918060 $T=23720 19910 0 0 $X=23500 $Y=19660
X156 82 M2_M1_CDNS_7656633918060 $T=23720 41110 0 0 $X=23500 $Y=40860
X157 83 M2_M1_CDNS_7656633918060 $T=26500 19910 0 0 $X=26280 $Y=19660
X158 84 M2_M1_CDNS_7656633918060 $T=26500 41110 0 0 $X=26280 $Y=40860
X159 85 M2_M1_CDNS_7656633918060 $T=36030 19910 0 0 $X=35810 $Y=19660
X160 86 M2_M1_CDNS_7656633918060 $T=36030 41110 0 0 $X=35810 $Y=40860
X161 87 M2_M1_CDNS_7656633918060 $T=44820 19910 0 0 $X=44600 $Y=19660
X162 88 M2_M1_CDNS_7656633918060 $T=44820 41110 0 0 $X=44600 $Y=40860
X163 89 M2_M1_CDNS_7656633918060 $T=50410 19910 0 0 $X=50190 $Y=19660
X164 90 M2_M1_CDNS_7656633918060 $T=50410 41110 0 0 $X=50190 $Y=40860
X165 91 M2_M1_CDNS_7656633918060 $T=53190 19910 0 0 $X=52970 $Y=19660
X166 92 M2_M1_CDNS_7656633918060 $T=53190 41110 0 0 $X=52970 $Y=40860
X167 78 M6_M5_CDNS_7656633918061 $T=9340 41110 0 0 $X=9120 $Y=40860
X168 79 M6_M5_CDNS_7656633918061 $T=18130 19910 0 0 $X=17910 $Y=19660
X169 80 M6_M5_CDNS_7656633918061 $T=18130 41110 0 0 $X=17910 $Y=40860
X170 81 M6_M5_CDNS_7656633918061 $T=23720 19910 0 0 $X=23500 $Y=19660
X171 82 M6_M5_CDNS_7656633918061 $T=23720 41110 0 0 $X=23500 $Y=40860
X172 83 M6_M5_CDNS_7656633918061 $T=26500 19910 0 0 $X=26280 $Y=19660
X173 84 M6_M5_CDNS_7656633918061 $T=26500 41110 0 0 $X=26280 $Y=40860
X174 85 M6_M5_CDNS_7656633918061 $T=36030 19910 0 0 $X=35810 $Y=19660
X175 86 M6_M5_CDNS_7656633918061 $T=36030 41110 0 0 $X=35810 $Y=40860
X176 87 M6_M5_CDNS_7656633918061 $T=44820 19910 0 0 $X=44600 $Y=19660
X177 88 M6_M5_CDNS_7656633918061 $T=44820 41110 0 0 $X=44600 $Y=40860
X178 89 M6_M5_CDNS_7656633918061 $T=50410 19910 0 0 $X=50190 $Y=19660
X179 90 M6_M5_CDNS_7656633918061 $T=50410 41110 0 0 $X=50190 $Y=40860
X180 91 M6_M5_CDNS_7656633918061 $T=53190 19910 0 0 $X=52970 $Y=19660
X181 92 M6_M5_CDNS_7656633918061 $T=53190 41110 0 0 $X=52970 $Y=40860
X182 6 1 4 3 78 107 183 AND $T=3670 43110 0 0 $X=4740 $Y=40010
X183 11 8 4 3 79 114 189 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X184 10 9 4 3 80 113 188 AND $T=12460 43110 0 0 $X=13530 $Y=40010
X185 17 14 4 3 81 120 195 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X186 16 15 4 3 82 119 194 AND $T=18050 43110 0 0 $X=19120 $Y=40010
X187 27 22 4 3 83 132 219 AND $T=32170 21910 1 180 $X=26920 $Y=18810
X188 26 23 4 3 84 131 218 AND $T=32170 43110 1 180 $X=26920 $Y=40010
X189 29 24 4 3 85 140 225 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X190 28 25 4 3 86 139 224 AND $T=30360 43110 0 0 $X=31430 $Y=40010
X191 35 32 4 3 87 146 233 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X192 34 33 4 3 88 145 232 AND $T=39150 43110 0 0 $X=40220 $Y=40010
X193 41 38 4 3 89 152 239 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X194 40 39 4 3 90 151 238 AND $T=44740 43110 0 0 $X=45810 $Y=40010
X195 45 48 4 3 91 159 246 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X196 44 49 4 3 92 158 245 AND $T=58860 43110 1 180 $X=53610 $Y=40010
X197 52 4 3 2 53 180 105 XOR $T=640 25900 1 0 $X=640 $Y=21200
X198 1 4 3 54 6 182 106 XOR $T=4740 40010 1 0 $X=4740 $Y=35310
X199 65 4 3 7 54 181 108 XOR $T=9740 25900 0 180 $X=6020 $Y=21200
X200 66 4 3 12 55 187 112 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X201 67 4 3 13 56 186 111 XOR $T=17180 25900 0 180 $X=13460 $Y=21200
X202 8 4 3 55 11 185 110 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X203 9 4 3 56 10 184 109 XOR $T=13530 40010 1 0 $X=13530 $Y=35310
X204 68 4 3 18 57 193 118 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X205 69 4 3 19 58 192 117 XOR $T=22760 25900 0 180 $X=19040 $Y=21200
X206 14 4 3 57 17 191 116 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X207 15 4 3 58 16 190 115 XOR $T=19120 40010 1 0 $X=19120 $Y=35310
X208 70 4 3 20 59 197 122 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X209 71 4 3 21 60 196 121 XOR $T=26810 25900 0 180 $X=23090 $Y=21200
X210 22 4 3 59 27 221 134 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X211 23 4 3 60 26 220 133 XOR $T=31140 40010 0 180 $X=27420 $Y=35310
X212 24 4 3 61 29 223 138 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X213 25 4 3 62 28 222 137 XOR $T=31430 40010 1 0 $X=31430 $Y=35310
X214 72 4 3 30 61 227 136 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X215 73 4 3 31 62 226 135 XOR $T=36470 25900 0 180 $X=32750 $Y=21200
X216 74 4 3 36 63 231 144 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X217 75 4 3 37 33 230 143 XOR $T=43890 25900 0 180 $X=40170 $Y=21200
X218 32 4 3 63 35 229 142 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X219 33 4 3 33 34 228 141 XOR $T=40220 40010 1 0 $X=40220 $Y=35310
X220 76 4 3 42 64 237 150 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X221 77 4 3 43 33 236 149 XOR $T=49450 25900 0 180 $X=45730 $Y=21200
X222 38 4 3 64 41 235 148 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X223 39 4 3 33 40 234 147 XOR $T=45810 40010 1 0 $X=45810 $Y=35310
X224 93 4 3 47 33 240 153 XOR $T=49650 25900 1 0 $X=49650 $Y=21200
X225 48 4 3 53 45 244 157 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X226 49 4 3 33 44 243 156 XOR $T=57790 40010 0 180 $X=54070 $Y=35310
X227 46 3 93 50 51 4 155 154 241 287
+ 288 242 HAdder $T=62720 27380 1 90 $X=53760 $Y=28180
X228 59 83 70 4 3 57 81 68 55 79
+ 66 94 5 95 96 101 102 103 104 257
+ 259 258 260 261 262 264 265 266 263 170
+ 171 174 175 173 176 177 172 178 179 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X229 60 84 71 4 3 58 82 69 56 80
+ 67 54 65 78 52 97 98 99 100 247
+ 249 248 250 251 252 254 255 256 253 160
+ 161 164 165 163 166 167 162 168 169 4bit_CLA_logic $T=26970 25900 1 180 $X=320 $Y=25900
X230 53 91 52 4 3 64 89 76 63 87
+ 74 61 72 85 70 127 128 129 130 277
+ 279 278 280 281 282 284 285 286 283 208
+ 209 212 213 211 214 215 210 216 217 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
X231 33 92 93 4 3 33 90 77 33 88
+ 75 62 73 86 71 123 124 125 126 267
+ 269 268 270 271 272 274 275 276 273 198
+ 199 202 203 201 204 205 200 206 207 4bit_CLA_logic $T=53660 25900 1 180 $X=27010 $Y=25900
M0 183 1 107 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5600 $Y=40350 $dt=0
M1 3 6 183 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=5810 $Y=40350 $dt=0
M2 78 107 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=8230 $Y=40340 $dt=0
M3 189 8 114 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=19150 $dt=0
M4 188 9 113 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14390 $Y=40350 $dt=0
M5 3 11 189 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=19150 $dt=0
M6 3 10 188 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=14600 $Y=40350 $dt=0
M7 79 114 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=19140 $dt=0
M8 80 113 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=17020 $Y=40340 $dt=0
M9 195 14 120 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=19150 $dt=0
M10 194 15 119 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=19980 $Y=40350 $dt=0
M11 3 17 195 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=19150 $dt=0
M12 3 16 194 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=20190 $Y=40350 $dt=0
M13 81 120 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=19140 $dt=0
M14 82 119 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=22610 $Y=40340 $dt=0
M15 3 132 83 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27520 $Y=19140 $dt=0
M16 3 131 84 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=27520 $Y=40340 $dt=0
M17 219 27 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29940 $Y=19150 $dt=0
M18 218 26 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=29940 $Y=40350 $dt=0
M19 132 22 219 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30150 $Y=19150 $dt=0
M20 131 23 218 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=30150 $Y=40350 $dt=0
M21 225 24 140 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=19150 $dt=0
M22 224 25 139 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32290 $Y=40350 $dt=0
M23 3 29 225 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=19150 $dt=0
M24 3 28 224 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=32500 $Y=40350 $dt=0
M25 85 140 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=19140 $dt=0
M26 86 139 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=34920 $Y=40340 $dt=0
M27 233 32 146 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=19150 $dt=0
M28 232 33 145 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41080 $Y=40350 $dt=0
M29 3 35 233 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=19150 $dt=0
M30 3 34 232 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=41290 $Y=40350 $dt=0
M31 87 146 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=19140 $dt=0
M32 88 145 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=43710 $Y=40340 $dt=0
M33 239 38 152 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=19150 $dt=0
M34 238 39 151 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46670 $Y=40350 $dt=0
M35 3 41 239 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=19150 $dt=0
M36 3 40 238 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=46880 $Y=40350 $dt=0
M37 89 152 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=19140 $dt=0
M38 90 151 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=49300 $Y=40340 $dt=0
M39 3 159 91 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=19140 $dt=0
M40 3 158 92 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=54210 $Y=40340 $dt=0
M41 246 45 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=19150 $dt=0
M42 245 44 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56630 $Y=40350 $dt=0
M43 159 48 246 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=19150 $dt=0
M44 158 49 245 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=56840 $Y=40350 $dt=0
M45 4 104 96 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M46 4 100 52 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=34270 $dt=1
M47 180 52 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=22000 $dt=1
M48 263 95 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M49 253 78 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=34270 $dt=1
M50 2 53 52 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=22000 $dt=1
M51 180 105 2 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=22000 $dt=1
M52 4 53 105 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=22000 $dt=1
M53 182 1 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=36110 $dt=1
M54 107 1 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=5600 $Y=41790 $dt=1
M55 4 6 107 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=6010 $Y=41790 $dt=1
M56 54 6 1 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=36110 $dt=1
M57 108 54 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=22000 $dt=1
M58 182 106 54 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=36110 $dt=1
M59 7 108 181 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=22000 $dt=1
M60 4 6 106 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=36110 $dt=1
M61 78 107 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=8230 $Y=41600 $dt=1
M62 65 54 7 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=22000 $dt=1
M63 4 65 181 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=22000 $dt=1
M64 112 55 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M65 111 56 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=115.144 scb=0.0588049 scc=0.0138331 $X=13880 $Y=22000 $dt=1
M66 185 8 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M67 184 9 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=36110 $dt=1
M68 114 8 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.29 scb=0.029437 scc=0.00332952 $X=14390 $Y=20590 $dt=1
M69 113 9 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=14390 $Y=41790 $dt=1
M70 4 11 114 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=28.0435 scb=0.0261338 scc=0.00329543 $X=14800 $Y=20590 $dt=1
M71 4 10 113 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=14800 $Y=41790 $dt=1
M72 12 112 187 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M73 13 111 186 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.854 scb=0.0354545 scc=0.011187 $X=14810 $Y=22000 $dt=1
M74 55 11 8 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M75 56 10 9 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=36110 $dt=1
M76 66 55 12 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M77 67 56 13 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=15740 $Y=22000 $dt=1
M78 185 110 55 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M79 184 109 56 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=36110 $dt=1
M80 4 66 187 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M81 4 67 186 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=16670 $Y=22000 $dt=1
M82 4 11 110 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M83 4 10 109 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=36110 $dt=1
M84 79 114 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=17020 $Y=20400 $dt=1
M85 80 113 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=17020 $Y=41600 $dt=1
M86 118 57 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M87 117 58 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=19460 $Y=22000 $dt=1
M88 191 14 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M89 190 15 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=36110 $dt=1
M90 120 14 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=19980 $Y=20590 $dt=1
M91 119 15 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=19980 $Y=41790 $dt=1
M92 18 118 193 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M93 4 17 120 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=20390 $Y=20590 $dt=1
M94 19 117 192 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=20390 $Y=22000 $dt=1
M95 4 16 119 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=20390 $Y=41790 $dt=1
M96 57 17 14 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M97 58 16 15 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=36110 $dt=1
M98 68 57 18 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M99 69 58 19 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=21320 $Y=22000 $dt=1
M100 191 116 57 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M101 190 115 58 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=36110 $dt=1
M102 4 68 193 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M103 4 69 192 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=22250 $Y=22000 $dt=1
M104 4 17 116 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M105 4 16 115 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=36110 $dt=1
M106 81 120 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=22610 $Y=20400 $dt=1
M107 82 119 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=22610 $Y=41600 $dt=1
M108 122 59 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M109 121 60 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=23510 $Y=22000 $dt=1
M110 20 122 197 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M111 21 121 196 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=24440 $Y=22000 $dt=1
M112 70 59 20 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M113 71 60 21 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=25370 $Y=22000 $dt=1
M114 4 70 197 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M115 4 71 196 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=26300 $Y=22000 $dt=1
M116 4 130 70 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M117 4 126 71 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=34270 $dt=1
M118 4 132 83 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=27520 $Y=20400 $dt=1
M119 4 131 84 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=27520 $Y=41600 $dt=1
M120 134 27 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M121 133 26 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=36110 $dt=1
M122 283 85 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M123 273 86 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=34270 $dt=1
M124 59 134 221 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M125 60 133 220 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=36110 $dt=1
M126 22 27 59 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M127 23 26 60 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=36110 $dt=1
M128 132 27 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=29740 $Y=20590 $dt=1
M129 131 26 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=29740 $Y=41790 $dt=1
M130 4 22 132 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=30150 $Y=20590 $dt=1
M131 4 23 131 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=30150 $Y=41790 $dt=1
M132 4 22 221 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M133 4 23 220 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=36110 $dt=1
M134 223 24 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M135 222 25 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=36110 $dt=1
M136 140 24 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32290 $Y=20590 $dt=1
M137 139 25 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32290 $Y=41790 $dt=1
M138 4 29 140 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32700 $Y=20590 $dt=1
M139 4 28 139 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32700 $Y=41790 $dt=1
M140 61 29 24 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M141 62 28 25 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=36110 $dt=1
M142 136 61 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M143 135 62 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=33170 $Y=22000 $dt=1
M144 223 138 61 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M145 222 137 62 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=36110 $dt=1
M146 30 136 227 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M147 31 135 226 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=34100 $Y=22000 $dt=1
M148 4 29 138 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M149 4 28 137 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=36110 $dt=1
M150 85 140 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=34920 $Y=20400 $dt=1
M151 86 139 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=34920 $Y=41600 $dt=1
M152 72 61 30 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M153 73 62 31 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35030 $Y=22000 $dt=1
M154 4 72 227 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M155 4 73 226 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35960 $Y=22000 $dt=1
M156 144 63 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M157 143 33 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=40590 $Y=22000 $dt=1
M158 229 32 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M159 228 33 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=36110 $dt=1
M160 146 32 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41080 $Y=20590 $dt=1
M161 145 33 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41080 $Y=41790 $dt=1
M162 4 35 146 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41490 $Y=20590 $dt=1
M163 4 34 145 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41490 $Y=41790 $dt=1
M164 36 144 231 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M165 37 143 230 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=41520 $Y=22000 $dt=1
M166 63 35 32 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M167 33 34 33 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=36110 $dt=1
M168 74 63 36 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M169 75 33 37 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=42450 $Y=22000 $dt=1
M170 229 142 63 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M171 228 141 33 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=36110 $dt=1
M172 4 74 231 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M173 4 75 230 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=43380 $Y=22000 $dt=1
M174 4 35 142 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M175 4 34 141 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=36110 $dt=1
M176 87 146 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=43710 $Y=20400 $dt=1
M177 88 145 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=43710 $Y=41600 $dt=1
M178 150 64 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M179 149 33 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=46150 $Y=22000 $dt=1
M180 235 38 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M181 234 39 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=36110 $dt=1
M182 152 38 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=46670 $Y=20590 $dt=1
M183 151 39 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=46670 $Y=41790 $dt=1
M184 42 150 237 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M185 4 41 152 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=47080 $Y=20590 $dt=1
M186 43 149 236 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=47080 $Y=22000 $dt=1
M187 4 40 151 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=47080 $Y=41790 $dt=1
M188 64 41 38 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M189 33 40 39 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=36110 $dt=1
M190 76 64 42 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=48010 $Y=800 $dt=1
M191 77 33 43 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48010 $Y=22000 $dt=1
M192 235 148 64 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M193 234 147 33 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=36110 $dt=1
M194 4 76 237 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=48940 $Y=800 $dt=1
M195 4 77 236 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48940 $Y=22000 $dt=1
M196 4 41 148 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M197 4 40 147 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=36110 $dt=1
M198 89 152 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=49300 $Y=20400 $dt=1
M199 90 151 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=49300 $Y=41600 $dt=1
M200 240 93 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=50070 $Y=22000 $dt=1
M201 47 33 93 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51000 $Y=22000 $dt=1
M202 240 153 47 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51930 $Y=22000 $dt=1
M203 4 33 153 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=52860 $Y=22000 $dt=1
M204 4 159 91 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=54210 $Y=20400 $dt=1
M205 4 158 92 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=54210 $Y=41600 $dt=1
M206 157 45 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M207 156 44 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=36110 $dt=1
M208 53 157 244 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M209 33 156 243 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=36110 $dt=1
M210 288 155 93 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=55830 $Y=32900 $dt=1
M211 4 154 288 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56040 $Y=32900 $dt=1
M212 48 45 53 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M213 49 44 33 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=36110 $dt=1
M214 159 45 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=29.0043 scb=0.0273456 scc=0.00330147 $X=56430 $Y=20590 $dt=1
M215 158 44 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=29.0043 scb=0.0273456 scc=0.00330147 $X=56430 $Y=41790 $dt=1
M216 4 48 159 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=33.5338 scb=0.0350848 scc=0.00355838 $X=56840 $Y=20590 $dt=1
M217 4 49 158 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=33.5338 scb=0.0350848 scc=0.00355838 $X=56840 $Y=41790 $dt=1
M218 4 154 287 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=56970 $Y=32900 $dt=1
M219 4 48 244 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M220 4 49 243 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=36110 $dt=1
M221 287 155 4 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57380 $Y=32900 $dt=1
M222 46 51 287 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=57790 $Y=32900 $dt=1
M223 287 50 46 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=58200 $Y=32900 $dt=1
M224 4 50 154 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=59130 $Y=32900 $dt=1
M225 4 51 155 4 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=60060 $Y=32900 $dt=1
.ends MAC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceProjectMAC                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceProjectMAC 198 197 196 195 194 193 192 191 190 200
+ 201 202 203 204 205 206 240 232 228 224
+ 222 216 212 235 231 227 223 221 215 211
+ 209 236 82 237 233 229 225 219 217 213
+ 208 238 234 230 226 220 218 214 210 207
+ 199 148 65 146 145 159 127 125 139 138
+ 140 147 75 74 64 149 80
** N=836 EP=67 FDC=2230
X0 1 M5_M4_CDNS_765663391800 $T=8680 96730 0 0 $X=8600 $Y=96600
X1 2 M5_M4_CDNS_765663391800 $T=17180 99960 0 0 $X=17100 $Y=99830
X2 3 M5_M4_CDNS_765663391800 $T=21730 98530 0 0 $X=21650 $Y=98400
X3 4 M5_M4_CDNS_765663391800 $T=25170 119910 0 0 $X=25090 $Y=119780
X4 5 M5_M4_CDNS_765663391800 $T=41900 93630 0 0 $X=41820 $Y=93500
X5 6 M5_M4_CDNS_765663391800 $T=42370 94030 0 0 $X=42290 $Y=93900
X6 7 M5_M4_CDNS_765663391800 $T=43570 92930 0 0 $X=43490 $Y=92800
X7 8 M5_M4_CDNS_765663391800 $T=43920 95730 0 0 $X=43840 $Y=95600
X8 9 M5_M4_CDNS_765663391800 $T=45720 98250 0 0 $X=45640 $Y=98120
X9 1 M5_M4_CDNS_765663391801 $T=8680 95430 0 0 $X=8550 $Y=95300
X10 10 M5_M4_CDNS_765663391801 $T=16520 72380 0 0 $X=16390 $Y=72250
X11 11 M5_M4_CDNS_765663391801 $T=19630 96730 0 0 $X=19500 $Y=96600
X12 8 M5_M4_CDNS_765663391801 $T=43920 101770 0 0 $X=43790 $Y=101640
X13 12 M4_M3_CDNS_765663391802 $T=2330 93930 0 0 $X=2200 $Y=93850
X14 13 M4_M3_CDNS_765663391802 $T=2680 98180 0 0 $X=2550 $Y=98100
X15 14 M4_M3_CDNS_765663391802 $T=6790 81230 0 0 $X=6660 $Y=81150
X16 15 M4_M3_CDNS_765663391802 $T=7630 101030 0 0 $X=7500 $Y=100950
X17 16 M4_M3_CDNS_765663391802 $T=8330 95080 0 0 $X=8200 $Y=95000
X18 1 M4_M3_CDNS_765663391802 $T=8680 95430 0 0 $X=8550 $Y=95350
X19 17 M4_M3_CDNS_765663391802 $T=9030 96030 0 0 $X=8900 $Y=95950
X20 8 M4_M3_CDNS_765663391802 $T=9730 95730 0 0 $X=9600 $Y=95650
X21 18 M4_M3_CDNS_765663391802 $T=10080 94280 0 0 $X=9950 $Y=94200
X22 7 M4_M3_CDNS_765663391802 $T=12540 92930 0 0 $X=12410 $Y=92850
X23 19 M4_M3_CDNS_765663391802 $T=15020 98900 0 0 $X=14890 $Y=98820
X24 5 M4_M3_CDNS_765663391802 $T=15890 93630 0 0 $X=15760 $Y=93550
X25 10 M4_M3_CDNS_765663391802 $T=16520 72380 0 0 $X=16390 $Y=72300
X26 20 M4_M3_CDNS_765663391802 $T=16890 86180 0 0 $X=16760 $Y=86100
X27 21 M4_M3_CDNS_765663391802 $T=17310 93230 0 0 $X=17180 $Y=93150
X28 12 M4_M3_CDNS_765663391802 $T=17310 93930 0 0 $X=17180 $Y=93850
X29 18 M4_M3_CDNS_765663391802 $T=17310 94280 0 0 $X=17180 $Y=94200
X30 22 M4_M3_CDNS_765663391802 $T=17310 94630 0 0 $X=17180 $Y=94550
X31 17 M4_M3_CDNS_765663391802 $T=17310 96030 0 0 $X=17180 $Y=95950
X32 23 M4_M3_CDNS_765663391802 $T=18510 99620 0 0 $X=18380 $Y=99540
X33 2 M4_M3_CDNS_765663391802 $T=18670 88620 0 0 $X=18540 $Y=88540
X34 24 M4_M3_CDNS_765663391802 $T=18930 99580 0 0 $X=18800 $Y=99500
X35 6 M4_M3_CDNS_765663391802 $T=19890 98480 0 0 $X=19760 $Y=98400
X36 23 M4_M3_CDNS_765663391802 $T=20680 81120 0 0 $X=20550 $Y=81040
X37 3 M4_M3_CDNS_765663391802 $T=22430 98530 0 0 $X=22300 $Y=98450
X38 25 M4_M3_CDNS_765663391802 $T=24660 97130 0 0 $X=24530 $Y=97050
X39 26 M4_M3_CDNS_765663391802 $T=25200 109890 0 0 $X=25070 $Y=109810
X40 27 M4_M3_CDNS_765663391802 $T=25740 97130 0 0 $X=25610 $Y=97050
X41 28 M4_M3_CDNS_765663391802 $T=25910 97830 0 0 $X=25780 $Y=97750
X42 29 M4_M3_CDNS_765663391802 $T=26000 113050 0 0 $X=25870 $Y=112970
X43 30 M4_M3_CDNS_765663391802 $T=27040 100570 0 0 $X=26910 $Y=100490
X44 31 M4_M3_CDNS_765663391802 $T=27410 101330 0 0 $X=27280 $Y=101250
X45 13 M4_M3_CDNS_765663391802 $T=29840 98180 0 0 $X=29710 $Y=98100
X46 19 M4_M3_CDNS_765663391802 $T=30510 93230 0 0 $X=30380 $Y=93150
X47 15 M4_M3_CDNS_765663391802 $T=31330 101030 0 0 $X=31200 $Y=100950
X48 32 M4_M3_CDNS_765663391802 $T=34650 79520 0 0 $X=34520 $Y=79440
X49 32 M4_M3_CDNS_765663391802 $T=34650 101010 0 0 $X=34520 $Y=100930
X50 33 M4_M3_CDNS_765663391802 $T=35310 99930 0 0 $X=35180 $Y=99850
X51 20 M4_M3_CDNS_765663391802 $T=37310 86180 0 0 $X=37180 $Y=86100
X52 34 M4_M3_CDNS_765663391802 $T=39310 85830 0 0 $X=39180 $Y=85750
X53 35 M4_M3_CDNS_765663391802 $T=40690 94330 0 0 $X=40560 $Y=94250
X54 11 M4_M3_CDNS_765663391802 $T=41190 96030 0 0 $X=41060 $Y=95950
X55 36 M4_M3_CDNS_765663391802 $T=42140 100630 0 0 $X=42010 $Y=100550
X56 24 M4_M3_CDNS_765663391802 $T=46090 99580 0 0 $X=45960 $Y=99500
X57 37 M4_M3_CDNS_765663391802 $T=46480 100160 0 0 $X=46350 $Y=100080
X58 38 M4_M3_CDNS_765663391802 $T=48490 98880 0 0 $X=48360 $Y=98800
X59 19 M5_M4_CDNS_765663391803 $T=15020 98900 0 0 $X=14890 $Y=98530
X60 10 M5_M4_CDNS_765663391803 $T=16520 91390 0 0 $X=16390 $Y=91020
X61 39 M5_M4_CDNS_765663391803 $T=16830 118300 0 0 $X=16700 $Y=117930
X62 40 M5_M4_CDNS_765663391803 $T=17570 117850 0 0 $X=17440 $Y=117480
X63 2 M5_M4_CDNS_765663391803 $T=18670 88620 0 0 $X=18540 $Y=88250
X64 40 M5_M4_CDNS_765663391803 $T=21030 80000 0 0 $X=20900 $Y=79630
X65 4 M5_M4_CDNS_765663391803 $T=25170 72590 0 0 $X=25040 $Y=72220
X66 32 M5_M4_CDNS_765663391803 $T=34650 79520 0 0 $X=34520 $Y=79150
X67 5 M5_M4_CDNS_765663391803 $T=41900 100280 0 0 $X=41770 $Y=99910
X68 6 M5_M4_CDNS_765663391803 $T=42370 100280 0 0 $X=42240 $Y=99910
X69 7 M5_M4_CDNS_765663391803 $T=43570 102040 0 0 $X=43440 $Y=101670
X70 21 M4_M3_CDNS_765663391804 $T=1900 93230 0 0 $X=1820 $Y=93100
X71 41 M4_M3_CDNS_765663391804 $T=3650 92530 0 0 $X=3570 $Y=92400
X72 42 M4_M3_CDNS_765663391804 $T=5880 82250 0 0 $X=5800 $Y=82120
X73 42 M4_M3_CDNS_765663391804 $T=5880 87300 0 0 $X=5800 $Y=87170
X74 43 M4_M3_CDNS_765663391804 $T=8380 96380 0 0 $X=8300 $Y=96250
X75 30 M4_M3_CDNS_765663391804 $T=10800 100570 0 0 $X=10720 $Y=100440
X76 44 M4_M3_CDNS_765663391804 $T=11190 74080 0 0 $X=11110 $Y=73950
X77 10 M4_M3_CDNS_765663391804 $T=16520 91390 0 0 $X=16440 $Y=91260
X78 2 M4_M3_CDNS_765663391804 $T=17180 100220 0 0 $X=17100 $Y=100090
X79 39 M4_M3_CDNS_765663391804 $T=21380 73000 0 0 $X=21300 $Y=72870
X80 45 M4_M3_CDNS_765663391804 $T=31390 100680 0 0 $X=31310 $Y=100550
X81 41 M4_M3_CDNS_765663391804 $T=41800 92530 0 0 $X=41720 $Y=92400
X82 9 M4_M3_CDNS_765663391804 $T=45720 98510 0 0 $X=45640 $Y=98380
X83 46 M4_M3_CDNS_765663391804 $T=47260 97130 0 0 $X=47180 $Y=97000
X84 31 M4_M3_CDNS_765663391804 $T=55100 101330 0 0 $X=55020 $Y=101200
X85 28 M4_M3_CDNS_765663391804 $T=59910 100550 0 0 $X=59830 $Y=100420
X86 22 M4_M3_CDNS_765663391805 $T=-390 94630 0 0 $X=-520 $Y=94260
X87 9 M4_M3_CDNS_765663391805 $T=3030 97480 0 0 $X=2900 $Y=97110
X88 47 M4_M3_CDNS_765663391805 $T=8310 71930 0 0 $X=8180 $Y=71560
X89 44 M4_M3_CDNS_765663391805 $T=11190 88980 0 0 $X=11060 $Y=88610
X90 29 M4_M3_CDNS_765663391805 $T=13830 111740 0 0 $X=13700 $Y=111370
X91 39 M4_M3_CDNS_765663391805 $T=16830 118300 0 0 $X=16700 $Y=117930
X92 38 M4_M3_CDNS_765663391805 $T=17310 98880 0 0 $X=17180 $Y=98510
X93 40 M4_M3_CDNS_765663391805 $T=17570 117850 0 0 $X=17440 $Y=117480
X94 33 M4_M3_CDNS_765663391805 $T=17580 99930 0 0 $X=17450 $Y=99560
X95 48 M4_M3_CDNS_765663391805 $T=18930 101770 0 0 $X=18800 $Y=101400
X96 35 M4_M3_CDNS_765663391805 $T=20130 103160 0 0 $X=20000 $Y=102790
X97 3 M4_M3_CDNS_765663391805 $T=20130 111380 0 0 $X=20000 $Y=111010
X98 49 M4_M3_CDNS_765663391805 $T=22690 99230 0 0 $X=22560 $Y=98860
X99 4 M4_M3_CDNS_765663391805 $T=25170 72590 0 0 $X=25040 $Y=72220
X100 43 M4_M3_CDNS_765663391805 $T=41190 100330 0 0 $X=41060 $Y=99960
X101 5 M4_M3_CDNS_765663391805 $T=41900 100280 0 0 $X=41770 $Y=99910
X102 6 M4_M3_CDNS_765663391805 $T=42370 100280 0 0 $X=42240 $Y=99910
X103 16 M4_M3_CDNS_765663391805 $T=42400 95080 0 0 $X=42270 $Y=94710
X104 37 M4_M3_CDNS_765663391805 $T=43230 100160 0 0 $X=43100 $Y=99790
X105 7 M4_M3_CDNS_765663391805 $T=43570 102040 0 0 $X=43440 $Y=101670
X106 34 M4_M3_CDNS_765663391805 $T=47850 88280 0 0 $X=47720 $Y=87910
X107 50 M3_M2_CDNS_765663391806 $T=1330 80160 0 0 $X=1250 $Y=80030
X108 50 M3_M2_CDNS_765663391806 $T=1330 104390 0 0 $X=1250 $Y=104260
X109 26 M3_M2_CDNS_765663391806 $T=2250 111070 0 0 $X=2170 $Y=110940
X110 26 M3_M2_CDNS_765663391806 $T=2250 112040 0 0 $X=2170 $Y=111910
X111 13 M3_M2_CDNS_765663391806 $T=2680 88600 0 0 $X=2600 $Y=88470
X112 9 M3_M2_CDNS_765663391806 $T=3030 97480 0 0 $X=2950 $Y=97350
X113 45 M3_M2_CDNS_765663391806 $T=4510 82980 0 0 $X=4430 $Y=82850
X114 51 M3_M2_CDNS_765663391806 $T=5010 87930 0 0 $X=4930 $Y=87800
X115 15 M3_M2_CDNS_765663391806 $T=6280 95080 0 0 $X=6200 $Y=94950
X116 16 M3_M2_CDNS_765663391806 $T=8330 95660 0 0 $X=8250 $Y=95530
X117 17 M3_M2_CDNS_765663391806 $T=9030 100590 0 0 $X=8950 $Y=100460
X118 8 M3_M2_CDNS_765663391806 $T=9730 98040 0 0 $X=9650 $Y=97910
X119 44 M3_M2_CDNS_765663391806 $T=11190 88980 0 0 $X=11110 $Y=88850
X120 52 M3_M2_CDNS_765663391806 $T=11410 96380 0 0 $X=11330 $Y=96250
X121 53 M3_M2_CDNS_765663391806 $T=11710 95430 0 0 $X=11630 $Y=95300
X122 53 M3_M2_CDNS_765663391806 $T=11710 97340 0 0 $X=11630 $Y=97210
X123 53 M3_M2_CDNS_765663391806 $T=11710 99520 0 0 $X=11630 $Y=99390
X124 7 M3_M2_CDNS_765663391806 $T=12540 94390 0 0 $X=12460 $Y=94260
X125 5 M3_M2_CDNS_765663391806 $T=15890 94270 0 0 $X=15810 $Y=94140
X126 39 M3_M2_CDNS_765663391806 $T=16830 118300 0 0 $X=16750 $Y=118170
X127 54 M3_M2_CDNS_765663391806 $T=16920 74000 0 0 $X=16840 $Y=73870
X128 1 M3_M2_CDNS_765663391806 $T=17100 96730 0 0 $X=17020 $Y=96600
X129 40 M3_M2_CDNS_765663391806 $T=17570 117850 0 0 $X=17490 $Y=117720
X130 33 M3_M2_CDNS_765663391806 $T=17580 99930 0 0 $X=17500 $Y=99800
X131 48 M3_M2_CDNS_765663391806 $T=18140 98310 0 0 $X=18060 $Y=98180
X132 48 M3_M2_CDNS_765663391806 $T=18140 99650 0 0 $X=18060 $Y=99520
X133 55 M3_M2_CDNS_765663391806 $T=21690 86530 0 0 $X=21610 $Y=86400
X134 34 M3_M2_CDNS_765663391806 $T=22040 85830 0 0 $X=21960 $Y=85700
X135 3 M3_M2_CDNS_765663391806 $T=22430 96730 0 0 $X=22350 $Y=96600
X136 49 M3_M2_CDNS_765663391806 $T=22690 99230 0 0 $X=22610 $Y=99100
X137 30 M3_M2_CDNS_765663391806 $T=27040 100380 0 0 $X=26960 $Y=100250
X138 31 M3_M2_CDNS_765663391806 $T=27410 98880 0 0 $X=27330 $Y=98750
X139 1 M3_M2_CDNS_765663391806 $T=29350 98980 0 0 $X=29270 $Y=98850
X140 19 M3_M2_CDNS_765663391806 $T=30510 93570 0 0 $X=30430 $Y=93440
X141 56 M3_M2_CDNS_765663391806 $T=31450 90030 0 0 $X=31370 $Y=89900
X142 42 M3_M2_CDNS_765663391806 $T=32290 87300 0 0 $X=32210 $Y=87170
X143 57 M3_M2_CDNS_765663391806 $T=35660 72840 0 0 $X=35580 $Y=72710
X144 58 M3_M2_CDNS_765663391806 $T=36230 101110 0 0 $X=36150 $Y=100980
X145 58 M3_M2_CDNS_765663391806 $T=36230 104400 0 0 $X=36150 $Y=104270
X146 59 M3_M2_CDNS_765663391806 $T=38790 101400 0 0 $X=38710 $Y=101270
X147 17 M3_M2_CDNS_765663391806 $T=39890 96030 0 0 $X=39810 $Y=95900
X148 35 M3_M2_CDNS_765663391806 $T=40690 96080 0 0 $X=40610 $Y=95950
X149 41 M3_M2_CDNS_765663391806 $T=41800 96430 0 0 $X=41720 $Y=96300
X150 16 M3_M2_CDNS_765663391806 $T=42400 95250 0 0 $X=42320 $Y=95120
X151 7 M3_M2_CDNS_765663391806 $T=43570 102040 0 0 $X=43490 $Y=101910
X152 8 M3_M2_CDNS_765663391806 $T=43920 101770 0 0 $X=43840 $Y=101640
X153 24 M3_M2_CDNS_765663391806 $T=46090 100580 0 0 $X=46010 $Y=100450
X154 60 M3_M2_CDNS_765663391806 $T=46110 91130 0 0 $X=46030 $Y=91000
X155 37 M3_M2_CDNS_765663391806 $T=46480 98530 0 0 $X=46400 $Y=98400
X156 61 M3_M2_CDNS_765663391806 $T=47390 96330 0 0 $X=47310 $Y=96200
X157 34 M3_M2_CDNS_765663391806 $T=47850 88280 0 0 $X=47770 $Y=88150
X158 38 M3_M2_CDNS_765663391806 $T=48490 99650 0 0 $X=48410 $Y=99520
X159 27 M3_M2_CDNS_765663391806 $T=49320 97160 0 0 $X=49240 $Y=97030
X160 31 M3_M2_CDNS_765663391806 $T=55100 100540 0 0 $X=55020 $Y=100410
X161 28 M3_M2_CDNS_765663391806 $T=59910 100810 0 0 $X=59830 $Y=100680
X162 37 M3_M2_CDNS_765663391806 $T=60410 97860 0 0 $X=60330 $Y=97730
X163 62 M3_M2_CDNS_765663391806 $T=60710 100630 0 0 $X=60630 $Y=100500
X164 19 M5_M4_CDNS_765663391807 $T=17730 94630 0 0 $X=17600 $Y=94550
X165 6 M5_M4_CDNS_765663391807 $T=19280 94030 0 0 $X=19150 $Y=93950
X166 6 M5_M4_CDNS_765663391807 $T=19280 98480 0 0 $X=19150 $Y=98400
X167 11 M5_M4_CDNS_765663391807 $T=19630 96030 0 0 $X=19500 $Y=95950
X168 23 M5_M4_CDNS_765663391807 $T=19980 81120 0 0 $X=19850 $Y=81040
X169 39 M5_M4_CDNS_765663391807 $T=21380 89430 0 0 $X=21250 $Y=89350
X170 3 M5_M4_CDNS_765663391807 $T=21730 111380 0 0 $X=21600 $Y=111300
X171 25 M5_M4_CDNS_765663391807 $T=24660 90430 0 0 $X=24530 $Y=90350
X172 19 M5_M4_CDNS_765663391807 $T=30510 94630 0 0 $X=30380 $Y=94550
X173 45 M5_M4_CDNS_765663391807 $T=31390 100230 0 0 $X=31260 $Y=100150
X174 36 M5_M4_CDNS_765663391807 $T=33310 100630 0 0 $X=33180 $Y=100550
X175 35 M5_M4_CDNS_765663391807 $T=40690 103160 0 0 $X=40560 $Y=103080
X176 43 M5_M4_CDNS_765663391807 $T=41190 96380 0 0 $X=41060 $Y=96300
X177 9 M5_M4_CDNS_765663391807 $T=45720 97480 0 0 $X=45590 $Y=97400
X178 63 M5_M4_CDNS_765663391808 $T=18230 111270 0 0 $X=18150 $Y=111020
X179 63 M5_M4_CDNS_765663391808 $T=20330 89330 0 0 $X=20250 $Y=89080
X180 2 M2_M1_CDNS_765663391809 $T=17180 111020 0 0 $X=17100 $Y=110770
X181 63 M2_M1_CDNS_765663391809 $T=18230 111270 0 0 $X=18150 $Y=111020
X182 48 M2_M1_CDNS_765663391809 $T=37450 101760 0 0 $X=37370 $Y=101510
X183 64 M4_M3_CDNS_7656633918010 $T=4820 42750 0 0 $X=4740 $Y=42500
X184 63 M4_M3_CDNS_7656633918010 $T=18230 111270 0 0 $X=18150 $Y=111020
X185 65 M4_M3_CDNS_7656633918010 $T=60960 21490 0 0 $X=60880 $Y=21240
X186 2 M3_M2_CDNS_7656633918011 $T=17180 111020 0 0 $X=17100 $Y=110770
X187 63 M3_M2_CDNS_7656633918011 $T=18230 111270 0 0 $X=18150 $Y=111020
X188 48 M3_M2_CDNS_7656633918011 $T=37450 101760 0 0 $X=37370 $Y=101510
X189 23 M5_M4_CDNS_7656633918012 $T=18510 99620 0 0 $X=18140 $Y=99490
X190 49 M5_M4_CDNS_7656633918012 $T=22690 99230 0 0 $X=22320 $Y=99100
X191 25 M5_M4_CDNS_7656633918012 $T=24660 97130 0 0 $X=24290 $Y=97000
X192 19 M5_M4_CDNS_7656633918012 $T=30510 93230 0 0 $X=30140 $Y=93100
X193 32 M5_M4_CDNS_7656633918012 $T=34650 101010 0 0 $X=34280 $Y=100880
X194 35 M5_M4_CDNS_7656633918012 $T=40690 94330 0 0 $X=40320 $Y=94200
X195 43 M5_M4_CDNS_7656633918012 $T=41190 100330 0 0 $X=40820 $Y=100200
X196 20 M4_M3_CDNS_7656633918013 $T=16890 88280 0 0 $X=16760 $Y=88150
X197 1 M4_M3_CDNS_7656633918013 $T=17100 96730 0 0 $X=16970 $Y=96600
X198 11 M4_M3_CDNS_7656633918013 $T=19630 96730 0 0 $X=19500 $Y=96600
X199 40 M4_M3_CDNS_7656633918013 $T=21030 80000 0 0 $X=20900 $Y=79870
X200 46 M4_M3_CDNS_7656633918013 $T=21270 96780 0 0 $X=21140 $Y=96650
X201 8 M4_M3_CDNS_7656633918013 $T=43920 101770 0 0 $X=43790 $Y=101640
X202 66 M3_M2_CDNS_7656633918014 $T=-700 73550 0 0 $X=-830 $Y=73180
X203 22 M3_M2_CDNS_7656633918014 $T=-390 94630 0 0 $X=-520 $Y=94260
X204 67 M3_M2_CDNS_7656633918014 $T=3160 89330 0 0 $X=3030 $Y=88960
X205 41 M3_M2_CDNS_7656633918014 $T=3650 90320 0 0 $X=3520 $Y=89950
X206 36 M3_M2_CDNS_7656633918014 $T=4000 89680 0 0 $X=3870 $Y=89310
X207 42 M3_M2_CDNS_7656633918014 $T=5880 81840 0 0 $X=5750 $Y=81470
X208 14 M3_M2_CDNS_7656633918014 $T=6580 110930 0 0 $X=6450 $Y=110560
X209 1 M3_M2_CDNS_7656633918014 $T=8790 112270 0 0 $X=8660 $Y=111900
X210 32 M3_M2_CDNS_7656633918014 $T=9930 79520 0 0 $X=9800 $Y=79150
X211 25 M3_M2_CDNS_7656633918014 $T=9950 90030 0 0 $X=9820 $Y=89660
X212 18 M3_M2_CDNS_7656633918014 $T=9950 111680 0 0 $X=9820 $Y=111310
X213 30 M3_M2_CDNS_7656633918014 $T=10800 97220 0 0 $X=10670 $Y=96850
X214 29 M3_M2_CDNS_7656633918014 $T=13830 111740 0 0 $X=13700 $Y=111370
X215 19 M3_M2_CDNS_7656633918014 $T=15160 111350 0 0 $X=15030 $Y=110980
X216 23 M3_M2_CDNS_7656633918014 $T=17880 118160 0 0 $X=17750 $Y=117790
X217 48 M3_M2_CDNS_7656633918014 $T=18930 101770 0 0 $X=18800 $Y=101400
X218 11 M3_M2_CDNS_7656633918014 $T=19630 96730 0 0 $X=19500 $Y=96360
X219 6 M3_M2_CDNS_7656633918014 $T=20550 98480 0 0 $X=20420 $Y=98110
X220 46 M3_M2_CDNS_7656633918014 $T=21270 96780 0 0 $X=21140 $Y=96410
X221 2 M3_M2_CDNS_7656633918014 $T=21290 88620 0 0 $X=21160 $Y=88250
X222 26 M3_M2_CDNS_7656633918014 $T=25200 101440 0 0 $X=25070 $Y=101070
X223 51 M3_M2_CDNS_7656633918014 $T=25520 88380 0 0 $X=25390 $Y=88010
X224 29 M3_M2_CDNS_7656633918014 $T=26000 101440 0 0 $X=25870 $Y=101070
X225 68 M3_M2_CDNS_7656633918014 $T=31890 98160 0 0 $X=31760 $Y=97790
X226 69 M3_M2_CDNS_7656633918014 $T=32630 79950 0 0 $X=32500 $Y=79580
X227 32 M3_M2_CDNS_7656633918014 $T=34650 101460 0 0 $X=34520 $Y=101090
X228 13 M3_M2_CDNS_7656633918014 $T=36630 99550 0 0 $X=36500 $Y=99180
X229 56 M3_M2_CDNS_7656633918014 $T=36860 88380 0 0 $X=36730 $Y=88010
X230 62 M3_M2_CDNS_7656633918014 $T=36940 96980 0 0 $X=36810 $Y=96610
X231 70 M3_M2_CDNS_7656633918014 $T=39070 97510 0 0 $X=38940 $Y=97140
X232 37 M3_M2_CDNS_7656633918014 $T=43230 100160 0 0 $X=43100 $Y=99790
X233 55 M3_M2_CDNS_7656633918014 $T=47850 80600 0 0 $X=47720 $Y=80230
X234 61 M3_M2_CDNS_7656633918014 $T=55310 88680 0 0 $X=55180 $Y=88310
X235 68 M3_M2_CDNS_7656633918014 $T=57720 100570 0 0 $X=57590 $Y=100200
X236 21 M3_M2_CDNS_7656633918017 $T=1900 111430 0 0 $X=1770 $Y=111350
X237 49 M3_M2_CDNS_7656633918017 $T=2490 82630 0 0 $X=2360 $Y=82550
X238 14 M3_M2_CDNS_7656633918017 $T=6580 95430 0 0 $X=6450 $Y=95350
X239 14 M3_M2_CDNS_7656633918017 $T=6790 89980 0 0 $X=6660 $Y=89900
X240 44 M3_M2_CDNS_7656633918017 $T=7280 95430 0 0 $X=7150 $Y=95350
X241 44 M3_M2_CDNS_7656633918017 $T=7280 107040 0 0 $X=7150 $Y=106960
X242 47 M3_M2_CDNS_7656633918017 $T=8310 71930 0 0 $X=8180 $Y=71850
X243 71 M3_M2_CDNS_7656633918017 $T=8960 90460 0 0 $X=8830 $Y=90380
X244 44 M3_M2_CDNS_7656633918017 $T=11190 71410 0 0 $X=11060 $Y=71330
X245 72 M3_M2_CDNS_7656633918017 $T=12880 91070 0 0 $X=12750 $Y=90990
X246 67 M3_M2_CDNS_7656633918017 $T=13310 89330 0 0 $X=13180 $Y=89250
X247 57 M3_M2_CDNS_7656633918017 $T=16450 81790 0 0 $X=16320 $Y=81710
X248 1 M3_M2_CDNS_7656633918017 $T=17100 95130 0 0 $X=16970 $Y=95050
X249 38 M3_M2_CDNS_7656633918017 $T=17310 98880 0 0 $X=17180 $Y=98800
X250 73 M3_M2_CDNS_7656633918017 $T=18260 80900 0 0 $X=18130 $Y=80820
X251 24 M3_M2_CDNS_7656633918017 $T=18930 99230 0 0 $X=18800 $Y=99150
X252 73 M3_M2_CDNS_7656633918017 $T=19940 80900 0 0 $X=19810 $Y=80820
X253 57 M3_M2_CDNS_7656633918017 $T=20310 81790 0 0 $X=20180 $Y=81710
X254 60 M3_M2_CDNS_7656633918017 $T=20540 91130 0 0 $X=20410 $Y=91050
X255 69 M3_M2_CDNS_7656633918017 $T=20680 80600 0 0 $X=20550 $Y=80520
X256 40 M3_M2_CDNS_7656633918017 $T=21030 80000 0 0 $X=20900 $Y=79920
X257 3 M3_M2_CDNS_7656633918017 $T=22430 95730 0 0 $X=22300 $Y=95650
X258 10 M3_M2_CDNS_7656633918017 $T=23880 90830 0 0 $X=23750 $Y=90750
X259 18 M3_M2_CDNS_7656633918017 $T=24330 94280 0 0 $X=24200 $Y=94200
X260 27 M3_M2_CDNS_7656633918017 $T=25170 97130 0 0 $X=25040 $Y=97050
X261 25 M3_M2_CDNS_7656633918017 $T=27010 96830 0 0 $X=26880 $Y=96750
X262 47 M3_M2_CDNS_7656633918017 $T=28680 91830 0 0 $X=28550 $Y=91750
X263 1 M3_M2_CDNS_7656633918017 $T=29350 95130 0 0 $X=29220 $Y=95050
X264 1 M3_M2_CDNS_7656633918017 $T=29350 101440 0 0 $X=29220 $Y=101360
X265 21 M3_M2_CDNS_7656633918017 $T=29800 93230 0 0 $X=29670 $Y=93150
X266 3 M3_M2_CDNS_7656633918017 $T=31030 95730 0 0 $X=30900 $Y=95650
X267 45 M3_M2_CDNS_7656633918017 $T=31170 100680 0 0 $X=31040 $Y=100600
X268 15 M3_M2_CDNS_7656633918017 $T=31610 101030 0 0 $X=31480 $Y=100950
X269 69 M3_M2_CDNS_7656633918017 $T=32630 80600 0 0 $X=32500 $Y=80520
X270 12 M3_M2_CDNS_7656633918017 $T=33720 93930 0 0 $X=33590 $Y=93850
X271 53 M3_M2_CDNS_7656633918017 $T=35430 95430 0 0 $X=35300 $Y=95350
X272 57 M3_M2_CDNS_7656633918017 $T=35660 81440 0 0 $X=35530 $Y=81360
X273 52 M3_M2_CDNS_7656633918017 $T=35830 96380 0 0 $X=35700 $Y=96300
X274 71 M3_M2_CDNS_7656633918017 $T=36510 90460 0 0 $X=36380 $Y=90380
X275 20 M3_M2_CDNS_7656633918017 $T=37310 88780 0 0 $X=37180 $Y=88700
X276 22 M3_M2_CDNS_7656633918017 $T=39490 94630 0 0 $X=39360 $Y=94550
X277 33 M3_M2_CDNS_7656633918017 $T=40290 99930 0 0 $X=40160 $Y=99850
X278 43 M3_M2_CDNS_7656633918017 $T=41190 100330 0 0 $X=41060 $Y=100250
X279 11 M3_M2_CDNS_7656633918017 $T=41450 96030 0 0 $X=41320 $Y=95950
X280 5 M3_M2_CDNS_7656633918017 $T=41900 100280 0 0 $X=41770 $Y=100200
X281 36 M3_M2_CDNS_7656633918017 $T=42400 100630 0 0 $X=42270 $Y=100550
X282 37 M3_M2_CDNS_7656633918017 $T=46480 97860 0 0 $X=46350 $Y=97780
X283 46 M3_M2_CDNS_7656633918017 $T=46830 97130 0 0 $X=46700 $Y=97050
X284 70 M3_M2_CDNS_7656633918017 $T=52950 97510 0 0 $X=52820 $Y=97430
X285 74 M5_M4_CDNS_7656633918018 $T=13070 42750 0 0 $X=12820 $Y=42670
X286 49 M5_M4_CDNS_7656633918018 $T=22690 82630 0 0 $X=22440 $Y=82550
X287 36 M5_M4_CDNS_7656633918018 $T=29310 89680 0 0 $X=29060 $Y=89600
X288 45 M5_M4_CDNS_7656633918018 $T=31390 82980 0 0 $X=31140 $Y=82900
X289 26 M4_M3_CDNS_7656633918019 $T=230 110810 0 0 $X=-20 $Y=110730
X290 75 M4_M3_CDNS_7656633918019 $T=18650 42750 0 0 $X=18400 $Y=42670
X291 49 M4_M3_CDNS_7656633918019 $T=22690 82630 0 0 $X=22440 $Y=82550
X292 47 M4_M3_CDNS_7656633918019 $T=28680 91830 0 0 $X=28430 $Y=91750
X293 36 M4_M3_CDNS_7656633918019 $T=29310 89680 0 0 $X=29060 $Y=89600
X294 45 M4_M3_CDNS_7656633918019 $T=31390 82980 0 0 $X=31140 $Y=82900
X295 66 M2_M1_CDNS_7656633918020 $T=-700 118270 0 0 $X=-780 $Y=118140
X296 76 M2_M1_CDNS_7656633918020 $T=-80 103430 0 0 $X=-160 $Y=103300
X297 66 M2_M1_CDNS_7656633918020 $T=1280 120900 0 0 $X=1200 $Y=120770
X298 13 M2_M1_CDNS_7656633918020 $T=1560 88600 0 0 $X=1480 $Y=88470
X299 26 M2_M1_CDNS_7656633918020 $T=2130 112300 0 0 $X=2050 $Y=112170
X300 49 M2_M1_CDNS_7656633918020 $T=2490 80510 0 0 $X=2410 $Y=80380
X301 9 M2_M1_CDNS_7656633918020 $T=2510 97480 0 0 $X=2430 $Y=97350
X302 77 M2_M1_CDNS_7656633918020 $T=2550 97970 0 0 $X=2470 $Y=97840
X303 51 M2_M1_CDNS_7656633918020 $T=2830 91250 0 0 $X=2750 $Y=91120
X304 76 M2_M1_CDNS_7656633918020 $T=2870 103430 0 0 $X=2790 $Y=103300
X305 78 M2_M1_CDNS_7656633918020 $T=3160 104950 0 0 $X=3080 $Y=104820
X306 79 M2_M1_CDNS_7656633918020 $T=3210 73020 0 0 $X=3130 $Y=72890
X307 80 M2_M1_CDNS_7656633918020 $T=3240 120790 0 0 $X=3160 $Y=120660
X308 78 M2_M1_CDNS_7656633918020 $T=3540 110950 0 0 $X=3460 $Y=110820
X309 41 M2_M1_CDNS_7656633918020 $T=3650 90320 0 0 $X=3570 $Y=90190
X310 45 M2_M1_CDNS_7656633918020 $T=4510 82170 0 0 $X=4430 $Y=82040
X311 69 M2_M1_CDNS_7656633918020 $T=5550 73490 0 0 $X=5470 $Y=73360
X312 80 M2_M1_CDNS_7656633918020 $T=6150 121230 0 0 $X=6070 $Y=121100
X313 81 M2_M1_CDNS_7656633918020 $T=6540 96610 0 0 $X=6460 $Y=96480
X314 81 M2_M1_CDNS_7656633918020 $T=6540 105070 0 0 $X=6460 $Y=104940
X315 14 M2_M1_CDNS_7656633918020 $T=6580 110930 0 0 $X=6500 $Y=110800
X316 73 M2_M1_CDNS_7656633918020 $T=6890 80900 0 0 $X=6810 $Y=80770
X317 16 M2_M1_CDNS_7656633918020 $T=8330 96510 0 0 $X=8250 $Y=96380
X318 43 M2_M1_CDNS_7656633918020 $T=8380 97010 0 0 $X=8300 $Y=96880
X319 69 M2_M1_CDNS_7656633918020 $T=8420 79410 0 0 $X=8340 $Y=79280
X320 1 M2_M1_CDNS_7656633918020 $T=8790 112270 0 0 $X=8710 $Y=112140
X321 82 M2_M1_CDNS_7656633918020 $T=8900 120860 0 0 $X=8820 $Y=120730
X322 8 M2_M1_CDNS_7656633918020 $T=9210 98040 0 0 $X=9130 $Y=97910
X323 25 M2_M1_CDNS_7656633918020 $T=9950 90030 0 0 $X=9870 $Y=89900
X324 18 M2_M1_CDNS_7656633918020 $T=9950 111680 0 0 $X=9870 $Y=111550
X325 44 M2_M1_CDNS_7656633918020 $T=10550 120910 0 0 $X=10470 $Y=120780
X326 52 M2_M1_CDNS_7656633918020 $T=11410 97340 0 0 $X=11330 $Y=97210
X327 52 M2_M1_CDNS_7656633918020 $T=11410 104450 0 0 $X=11330 $Y=104320
X328 82 M2_M1_CDNS_7656633918020 $T=11820 121150 0 0 $X=11740 $Y=121020
X329 7 M2_M1_CDNS_7656633918020 $T=12540 96660 0 0 $X=12460 $Y=96530
X330 72 M2_M1_CDNS_7656633918020 $T=12880 82460 0 0 $X=12800 $Y=82330
X331 39 M2_M1_CDNS_7656633918020 $T=13220 120920 0 0 $X=13140 $Y=120790
X332 44 M2_M1_CDNS_7656633918020 $T=13830 71410 0 0 $X=13750 $Y=71280
X333 29 M2_M1_CDNS_7656633918020 $T=13830 111740 0 0 $X=13750 $Y=111610
X334 80 M2_M1_CDNS_7656633918020 $T=14580 120890 0 0 $X=14500 $Y=120760
X335 80 M2_M1_CDNS_7656633918020 $T=15410 120950 0 0 $X=15330 $Y=120820
X336 83 M2_M1_CDNS_7656633918020 $T=15840 90790 0 0 $X=15760 $Y=90660
X337 5 M2_M1_CDNS_7656633918020 $T=15890 96510 0 0 $X=15810 $Y=96380
X338 40 M2_M1_CDNS_7656633918020 $T=16200 120910 0 0 $X=16120 $Y=120780
X339 84 M2_M1_CDNS_7656633918020 $T=16370 79450 0 0 $X=16290 $Y=79320
X340 84 M2_M1_CDNS_7656633918020 $T=17860 71590 0 0 $X=17780 $Y=71460
X341 84 M2_M1_CDNS_7656633918020 $T=17860 75760 0 0 $X=17780 $Y=75630
X342 23 M2_M1_CDNS_7656633918020 $T=18910 120910 0 0 $X=18830 $Y=120780
X343 11 M2_M1_CDNS_7656633918020 $T=19630 96660 0 0 $X=19550 $Y=96530
X344 3 M2_M1_CDNS_7656633918020 $T=20130 111380 0 0 $X=20050 $Y=111250
X345 82 M2_M1_CDNS_7656633918020 $T=20250 120910 0 0 $X=20170 $Y=120780
X346 60 M2_M1_CDNS_7656633918020 $T=20540 90800 0 0 $X=20460 $Y=90670
X347 6 M2_M1_CDNS_7656633918020 $T=20550 98480 0 0 $X=20470 $Y=98350
X348 55 M2_M1_CDNS_7656633918020 $T=20620 91480 0 0 $X=20540 $Y=91350
X349 46 M2_M1_CDNS_7656633918020 $T=21270 96660 0 0 $X=21190 $Y=96530
X350 2 M2_M1_CDNS_7656633918020 $T=21290 88620 0 0 $X=21210 $Y=88490
X351 39 M2_M1_CDNS_7656633918020 $T=21380 72640 0 0 $X=21300 $Y=72510
X352 4 M2_M1_CDNS_7656633918020 $T=21890 120910 0 0 $X=21810 $Y=120780
X353 34 M2_M1_CDNS_7656633918020 $T=22040 88140 0 0 $X=21960 $Y=88010
X354 85 M2_M1_CDNS_7656633918020 $T=22380 111680 0 0 $X=22300 $Y=111550
X355 58 M2_M1_CDNS_7656633918020 $T=22680 104400 0 0 $X=22600 $Y=104270
X356 82 M2_M1_CDNS_7656633918020 $T=23170 121220 0 0 $X=23090 $Y=121090
X357 10 M2_M1_CDNS_7656633918020 $T=23880 96990 0 0 $X=23800 $Y=96860
X358 18 M2_M1_CDNS_7656633918020 $T=24330 96980 0 0 $X=24250 $Y=96850
X359 4 M2_M1_CDNS_7656633918020 $T=25170 72590 0 0 $X=25090 $Y=72460
X360 26 M2_M1_CDNS_7656633918020 $T=25200 101440 0 0 $X=25120 $Y=101310
X361 51 M2_M1_CDNS_7656633918020 $T=25520 88380 0 0 $X=25440 $Y=88250
X362 86 M2_M1_CDNS_7656633918020 $T=25910 81790 0 0 $X=25830 $Y=81660
X363 29 M2_M1_CDNS_7656633918020 $T=26000 101440 0 0 $X=25920 $Y=101310
X364 31 M2_M1_CDNS_7656633918020 $T=26330 98880 0 0 $X=26250 $Y=98750
X365 85 M2_M1_CDNS_7656633918020 $T=26400 101440 0 0 $X=26320 $Y=101310
X366 49 M2_M1_CDNS_7656633918020 $T=26660 100640 0 0 $X=26580 $Y=100510
X367 25 M2_M1_CDNS_7656633918020 $T=27220 96830 0 0 $X=27140 $Y=96700
X368 83 M2_M1_CDNS_7656633918020 $T=27600 97880 0 0 $X=27520 $Y=97750
X369 47 M2_M1_CDNS_7656633918020 $T=28680 99330 0 0 $X=28600 $Y=99200
X370 21 M2_M1_CDNS_7656633918020 $T=29800 99700 0 0 $X=29720 $Y=99570
X371 87 M2_M1_CDNS_7656633918020 $T=30580 79400 0 0 $X=30500 $Y=79270
X372 3 M2_M1_CDNS_7656633918020 $T=31030 99380 0 0 $X=30950 $Y=99250
X373 88 M2_M1_CDNS_7656633918020 $T=31470 98510 0 0 $X=31390 $Y=98380
X374 15 M2_M1_CDNS_7656633918020 $T=31820 101030 0 0 $X=31740 $Y=100900
X375 89 M2_M1_CDNS_7656633918020 $T=31890 89330 0 0 $X=31810 $Y=89200
X376 42 M2_M1_CDNS_7656633918020 $T=32290 88570 0 0 $X=32210 $Y=88440
X377 69 M2_M1_CDNS_7656633918020 $T=32630 79950 0 0 $X=32550 $Y=79820
X378 12 M2_M1_CDNS_7656633918020 $T=33720 96520 0 0 $X=33640 $Y=96390
X379 57 M2_M1_CDNS_7656633918020 $T=35660 72580 0 0 $X=35580 $Y=72450
X380 58 M2_M1_CDNS_7656633918020 $T=36230 100850 0 0 $X=36150 $Y=100720
X381 71 M2_M1_CDNS_7656633918020 $T=36510 90170 0 0 $X=36430 $Y=90040
X382 13 M2_M1_CDNS_7656633918020 $T=36630 99550 0 0 $X=36550 $Y=99420
X383 56 M2_M1_CDNS_7656633918020 $T=36860 88380 0 0 $X=36780 $Y=88250
X384 62 M2_M1_CDNS_7656633918020 $T=36940 96980 0 0 $X=36860 $Y=96850
X385 30 M2_M1_CDNS_7656633918020 $T=37020 100380 0 0 $X=36940 $Y=100250
X386 59 M2_M1_CDNS_7656633918020 $T=38790 100280 0 0 $X=38710 $Y=100150
X387 70 M2_M1_CDNS_7656633918020 $T=39070 97510 0 0 $X=38990 $Y=97380
X388 22 M2_M1_CDNS_7656633918020 $T=39490 97070 0 0 $X=39410 $Y=96940
X389 90 M2_M1_CDNS_7656633918020 $T=39570 89330 0 0 $X=39490 $Y=89200
X390 17 M2_M1_CDNS_7656633918020 $T=39890 96740 0 0 $X=39810 $Y=96610
X391 33 M2_M1_CDNS_7656633918020 $T=40290 100140 0 0 $X=40210 $Y=100010
X392 35 M2_M1_CDNS_7656633918020 $T=40690 96700 0 0 $X=40610 $Y=96570
X393 91 M2_M1_CDNS_7656633918020 $T=40910 81680 0 0 $X=40830 $Y=81550
X394 92 M2_M1_CDNS_7656633918020 $T=40910 90200 0 0 $X=40830 $Y=90070
X395 41 M2_M1_CDNS_7656633918020 $T=41090 98880 0 0 $X=41010 $Y=98750
X396 43 M2_M1_CDNS_7656633918020 $T=41490 100330 0 0 $X=41410 $Y=100200
X397 5 M2_M1_CDNS_7656633918020 $T=41900 100920 0 0 $X=41820 $Y=100790
X398 11 M2_M1_CDNS_7656633918020 $T=42280 101440 0 0 $X=42200 $Y=101310
X399 6 M2_M1_CDNS_7656633918020 $T=42370 100280 0 0 $X=42290 $Y=100150
X400 93 M2_M1_CDNS_7656633918020 $T=43230 81310 0 0 $X=43150 $Y=81180
X401 37 M2_M1_CDNS_7656633918020 $T=43230 100160 0 0 $X=43150 $Y=100030
X402 94 M2_M1_CDNS_7656633918020 $T=43250 63930 0 0 $X=43170 $Y=63800
X403 7 M2_M1_CDNS_7656633918020 $T=43570 101180 0 0 $X=43490 $Y=101050
X404 20 M2_M1_CDNS_7656633918020 $T=43970 88780 0 0 $X=43890 $Y=88650
X405 95 M2_M1_CDNS_7656633918020 $T=43970 97220 0 0 $X=43890 $Y=97090
X406 36 M2_M1_CDNS_7656633918020 $T=45790 100630 0 0 $X=45710 $Y=100500
X407 24 M2_M1_CDNS_7656633918020 $T=46570 101430 0 0 $X=46490 $Y=101300
X408 46 M2_M1_CDNS_7656633918020 $T=46830 100430 0 0 $X=46750 $Y=100300
X409 61 M2_M1_CDNS_7656633918020 $T=47390 100770 0 0 $X=47310 $Y=100640
X410 96 M2_M1_CDNS_7656633918020 $T=47850 97220 0 0 $X=47770 $Y=97090
X411 97 M2_M1_CDNS_7656633918020 $T=47870 72330 0 0 $X=47790 $Y=72200
X412 98 M2_M1_CDNS_7656633918020 $T=48520 63930 0 0 $X=48440 $Y=63800
X413 91 M2_M1_CDNS_7656633918020 $T=48590 81680 0 0 $X=48510 $Y=81550
X414 99 M2_M1_CDNS_7656633918020 $T=48600 97620 0 0 $X=48520 $Y=97490
X415 100 M2_M1_CDNS_7656633918020 $T=50910 71610 0 0 $X=50830 $Y=71480
X416 101 M2_M1_CDNS_7656633918020 $T=50910 82090 0 0 $X=50830 $Y=81960
X417 102 M2_M1_CDNS_7656633918020 $T=50910 88980 0 0 $X=50830 $Y=88850
X418 103 M2_M1_CDNS_7656633918020 $T=50910 100060 0 0 $X=50830 $Y=99930
X419 59 M2_M1_CDNS_7656633918020 $T=51300 101460 0 0 $X=51220 $Y=101330
X420 95 M2_M1_CDNS_7656633918020 $T=51700 99890 0 0 $X=51620 $Y=99760
X421 96 M2_M1_CDNS_7656633918020 $T=52090 101040 0 0 $X=52010 $Y=100910
X422 104 M2_M1_CDNS_7656633918020 $T=54160 79510 0 0 $X=54080 $Y=79380
X423 104 M2_M1_CDNS_7656633918020 $T=54160 81970 0 0 $X=54080 $Y=81840
X424 9 M2_M1_CDNS_7656633918020 $T=54300 101520 0 0 $X=54220 $Y=101390
X425 105 M2_M1_CDNS_7656633918020 $T=54500 97910 0 0 $X=54420 $Y=97780
X426 102 M2_M1_CDNS_7656633918020 $T=54570 88980 0 0 $X=54490 $Y=88850
X427 31 M2_M1_CDNS_7656633918020 $T=55100 100280 0 0 $X=55020 $Y=100150
X428 61 M2_M1_CDNS_7656633918020 $T=55310 88680 0 0 $X=55230 $Y=88550
X429 70 M2_M1_CDNS_7656633918020 $T=55910 99800 0 0 $X=55830 $Y=99670
X430 105 M2_M1_CDNS_7656633918020 $T=56300 100030 0 0 $X=56220 $Y=99900
X431 106 M2_M1_CDNS_7656633918020 $T=56420 80850 0 0 $X=56340 $Y=80720
X432 107 M2_M1_CDNS_7656633918020 $T=56700 100940 0 0 $X=56620 $Y=100810
X433 108 M2_M1_CDNS_7656633918020 $T=57090 99720 0 0 $X=57010 $Y=99590
X434 109 M2_M1_CDNS_7656633918020 $T=59200 71290 0 0 $X=59120 $Y=71160
X435 110 M2_M1_CDNS_7656633918020 $T=59200 98490 0 0 $X=59120 $Y=98360
X436 111 M2_M1_CDNS_7656633918020 $T=59210 88110 0 0 $X=59130 $Y=87980
X437 28 M2_M1_CDNS_7656633918020 $T=59910 101100 0 0 $X=59830 $Y=100970
X438 62 M2_M1_CDNS_7656633918020 $T=60710 100970 0 0 $X=60630 $Y=100840
X439 37 M2_M1_CDNS_7656633918020 $T=61110 100660 0 0 $X=61030 $Y=100530
X440 43 M3_M2_CDNS_7656633918021 $T=8380 97010 0 0 $X=8010 $Y=96880
X441 10 M3_M2_CDNS_7656633918021 $T=16310 72380 0 0 $X=15940 $Y=72250
X442 20 M3_M2_CDNS_7656633918021 $T=16890 88280 0 0 $X=16520 $Y=88150
X443 54 M3_M2_CDNS_7656633918021 $T=20550 72330 0 0 $X=20180 $Y=72200
X444 4 M3_M2_CDNS_7656633918021 $T=25170 72590 0 0 $X=24800 $Y=72460
X445 23 M3_M2_CDNS_7656633918021 $T=25170 80000 0 0 $X=24800 $Y=79870
X446 66 M2_M1_CDNS_7656633918023 $T=-700 73550 0 0 $X=-830 $Y=73470
X447 22 M2_M1_CDNS_7656633918023 $T=-390 94630 0 0 $X=-520 $Y=94550
X448 22 M2_M1_CDNS_7656633918023 $T=-390 111110 0 0 $X=-520 $Y=111030
X449 76 M2_M1_CDNS_7656633918023 $T=-80 65150 0 0 $X=-210 $Y=65070
X450 112 M2_M1_CDNS_7656633918023 $T=230 71260 0 0 $X=100 $Y=71180
X451 22 M2_M1_CDNS_7656633918023 $T=1380 111110 0 0 $X=1250 $Y=111030
X452 47 M2_M1_CDNS_7656633918023 $T=2510 71930 0 0 $X=2380 $Y=71850
X453 50 M2_M1_CDNS_7656633918023 $T=2550 104900 0 0 $X=2420 $Y=104820
X454 21 M2_M1_CDNS_7656633918023 $T=2620 111430 0 0 $X=2490 $Y=111350
X455 76 M2_M1_CDNS_7656633918023 $T=3160 65150 0 0 $X=3030 $Y=65070
X456 67 M2_M1_CDNS_7656633918023 $T=3160 89330 0 0 $X=3030 $Y=89250
X457 36 M2_M1_CDNS_7656633918023 $T=4000 89680 0 0 $X=3870 $Y=89600
X458 10 M2_M1_CDNS_7656633918023 $T=4110 72380 0 0 $X=3980 $Y=72300
X459 38 M2_M1_CDNS_7656633918023 $T=4200 96710 0 0 $X=4070 $Y=96630
X460 42 M2_M1_CDNS_7656633918023 $T=5880 81840 0 0 $X=5750 $Y=81760
X461 113 M2_M1_CDNS_7656633918023 $T=5910 103750 0 0 $X=5780 $Y=103670
X462 112 M2_M1_CDNS_7656633918023 $T=6530 71260 0 0 $X=6400 $Y=71180
X463 81 M2_M1_CDNS_7656633918023 $T=6540 82200 0 0 $X=6410 $Y=82120
X464 71 M2_M1_CDNS_7656633918023 $T=7650 90460 0 0 $X=7520 $Y=90380
X465 69 M2_M1_CDNS_7656633918023 $T=8420 80300 0 0 $X=8290 $Y=80220
X466 15 M2_M1_CDNS_7656633918023 $T=8790 89080 0 0 $X=8660 $Y=89000
X467 17 M2_M1_CDNS_7656633918023 $T=8790 100590 0 0 $X=8660 $Y=100510
X468 57 M2_M1_CDNS_7656633918023 $T=9230 81790 0 0 $X=9100 $Y=81710
X469 66 M2_M1_CDNS_7656633918023 $T=9710 73550 0 0 $X=9580 $Y=73470
X470 32 M2_M1_CDNS_7656633918023 $T=9930 79520 0 0 $X=9800 $Y=79440
X471 53 M2_M1_CDNS_7656633918023 $T=9950 99520 0 0 $X=9820 $Y=99440
X472 114 M2_M1_CDNS_7656633918023 $T=10020 72080 0 0 $X=9890 $Y=72000
X473 30 M2_M1_CDNS_7656633918023 $T=10800 97220 0 0 $X=10670 $Y=97140
X474 52 M2_M1_CDNS_7656633918023 $T=13830 104450 0 0 $X=13700 $Y=104370
X475 50 M2_M1_CDNS_7656633918023 $T=13850 79870 0 0 $X=13720 $Y=79790
X476 54 M2_M1_CDNS_7656633918023 $T=13890 74000 0 0 $X=13760 $Y=73920
X477 115 M2_M1_CDNS_7656633918023 $T=13890 82600 0 0 $X=13760 $Y=82520
X478 114 M2_M1_CDNS_7656633918023 $T=14570 72080 0 0 $X=14440 $Y=72000
X479 24 M2_M1_CDNS_7656633918023 $T=14570 99230 0 0 $X=14440 $Y=99150
X480 33 M2_M1_CDNS_7656633918023 $T=14990 99930 0 0 $X=14860 $Y=99850
X481 19 M2_M1_CDNS_7656633918023 $T=15160 111350 0 0 $X=15030 $Y=111270
X482 48 M2_M1_CDNS_7656633918023 $T=15540 97390 0 0 $X=15410 $Y=97310
X483 20 M2_M1_CDNS_7656633918023 $T=16890 88280 0 0 $X=16760 $Y=88200
X484 116 M2_M1_CDNS_7656633918023 $T=18230 72030 0 0 $X=18100 $Y=71950
X485 14 M2_M1_CDNS_7656633918023 $T=18260 81230 0 0 $X=18130 $Y=81150
X486 86 M2_M1_CDNS_7656633918023 $T=18960 81490 0 0 $X=18830 $Y=81410
X487 67 M2_M1_CDNS_7656633918023 $T=20130 89330 0 0 $X=20000 $Y=89250
X488 35 M2_M1_CDNS_7656633918023 $T=20130 103160 0 0 $X=20000 $Y=103080
X489 54 M2_M1_CDNS_7656633918023 $T=20550 72330 0 0 $X=20420 $Y=72250
X490 86 M2_M1_CDNS_7656633918023 $T=22920 81490 0 0 $X=22790 $Y=81410
X491 86 M2_M1_CDNS_7656633918023 $T=22920 82090 0 0 $X=22790 $Y=82010
X492 113 M2_M1_CDNS_7656633918023 $T=24390 101500 0 0 $X=24260 $Y=101420
X493 23 M2_M1_CDNS_7656633918023 $T=25170 80000 0 0 $X=25040 $Y=79920
X494 27 M2_M1_CDNS_7656633918023 $T=25170 97280 0 0 $X=25040 $Y=97200
X495 117 M2_M1_CDNS_7656633918023 $T=25890 64850 0 0 $X=25760 $Y=64770
X496 116 M2_M1_CDNS_7656633918023 $T=25910 72030 0 0 $X=25780 $Y=71950
X497 28 M2_M1_CDNS_7656633918023 $T=25910 97510 0 0 $X=25780 $Y=97430
X498 118 M2_M1_CDNS_7656633918023 $T=28230 72030 0 0 $X=28100 $Y=71950
X499 87 M2_M1_CDNS_7656633918023 $T=28230 79400 0 0 $X=28100 $Y=79320
X500 89 M2_M1_CDNS_7656633918023 $T=28230 89330 0 0 $X=28100 $Y=89250
X501 119 M2_M1_CDNS_7656633918023 $T=29570 73370 0 0 $X=29440 $Y=73290
X502 120 M2_M1_CDNS_7656633918023 $T=29570 81860 0 0 $X=29440 $Y=81780
X503 56 M2_M1_CDNS_7656633918023 $T=29570 90030 0 0 $X=29440 $Y=89950
X504 19 M2_M1_CDNS_7656633918023 $T=30510 99330 0 0 $X=30380 $Y=99250
X505 45 M2_M1_CDNS_7656633918023 $T=31430 100680 0 0 $X=31300 $Y=100600
X506 118 M2_M1_CDNS_7656633918023 $T=31890 72030 0 0 $X=31760 $Y=71950
X507 68 M2_M1_CDNS_7656633918023 $T=31890 98160 0 0 $X=31760 $Y=98080
X508 79 M2_M1_CDNS_7656633918023 $T=32630 73020 0 0 $X=32500 $Y=72940
X509 103 M2_M1_CDNS_7656633918023 $T=32630 97180 0 0 $X=32500 $Y=97100
X510 32 M2_M1_CDNS_7656633918023 $T=34650 101460 0 0 $X=34520 $Y=101380
X511 119 M2_M1_CDNS_7656633918023 $T=35300 73370 0 0 $X=35170 $Y=73290
X512 53 M2_M1_CDNS_7656633918023 $T=35430 96890 0 0 $X=35300 $Y=96810
X513 52 M2_M1_CDNS_7656633918023 $T=35830 97110 0 0 $X=35700 $Y=97030
X514 73 M2_M1_CDNS_7656633918023 $T=36510 80900 0 0 $X=36380 $Y=80820
X515 120 M2_M1_CDNS_7656633918023 $T=37250 81860 0 0 $X=37120 $Y=81780
X516 121 M2_M1_CDNS_7656633918023 $T=39570 72030 0 0 $X=39440 $Y=71950
X517 93 M2_M1_CDNS_7656633918023 $T=39570 81310 0 0 $X=39440 $Y=81230
X518 97 M2_M1_CDNS_7656633918023 $T=40910 72330 0 0 $X=40780 $Y=72250
X519 88 M2_M1_CDNS_7656633918023 $T=41210 98510 0 0 $X=41080 $Y=98430
X520 121 M2_M1_CDNS_7656633918023 $T=43230 72030 0 0 $X=43100 $Y=71950
X521 90 M2_M1_CDNS_7656633918023 $T=43230 89330 0 0 $X=43100 $Y=89250
X522 8 M2_M1_CDNS_7656633918023 $T=43920 101480 0 0 $X=43790 $Y=101400
X523 84 M2_M1_CDNS_7656633918023 $T=43970 71590 0 0 $X=43840 $Y=71510
X524 115 M2_M1_CDNS_7656633918023 $T=43970 80300 0 0 $X=43840 $Y=80220
X525 95 M2_M1_CDNS_7656633918023 $T=43970 98920 0 0 $X=43840 $Y=98840
X526 16 M2_M1_CDNS_7656633918023 $T=44250 100050 0 0 $X=44120 $Y=99970
X527 60 M2_M1_CDNS_7656633918023 $T=46480 100080 0 0 $X=46350 $Y=100000
X528 55 M2_M1_CDNS_7656633918023 $T=47850 80600 0 0 $X=47720 $Y=80520
X529 34 M2_M1_CDNS_7656633918023 $T=47850 88570 0 0 $X=47720 $Y=88490
X530 122 M2_M1_CDNS_7656633918023 $T=47980 64630 0 0 $X=47850 $Y=64550
X531 92 M2_M1_CDNS_7656633918023 $T=48590 90200 0 0 $X=48460 $Y=90120
X532 99 M2_M1_CDNS_7656633918023 $T=48600 99300 0 0 $X=48470 $Y=99220
X533 27 M2_M1_CDNS_7656633918023 $T=49320 99840 0 0 $X=49190 $Y=99760
X534 107 M2_M1_CDNS_7656633918023 $T=51270 96980 0 0 $X=51140 $Y=96900
X535 95 M2_M1_CDNS_7656633918023 $T=51700 98920 0 0 $X=51570 $Y=98840
X536 101 M2_M1_CDNS_7656633918023 $T=51940 82090 0 0 $X=51810 $Y=82010
X537 108 M2_M1_CDNS_7656633918023 $T=53770 97030 0 0 $X=53640 $Y=96950
X538 123 M2_M1_CDNS_7656633918023 $T=54180 98860 0 0 $X=54050 $Y=98780
X539 123 M2_M1_CDNS_7656633918023 $T=54180 100120 0 0 $X=54050 $Y=100040
X540 124 M2_M1_CDNS_7656633918023 $T=55000 97030 0 0 $X=54870 $Y=96950
X541 109 M2_M1_CDNS_7656633918023 $T=55250 73700 0 0 $X=55120 $Y=73620
X542 100 M2_M1_CDNS_7656633918023 $T=55290 71610 0 0 $X=55160 $Y=71530
X543 68 M2_M1_CDNS_7656633918023 $T=57720 100570 0 0 $X=57590 $Y=100490
X544 110 M2_M1_CDNS_7656633918023 $T=58070 101400 0 0 $X=57940 $Y=101320
X545 106 M2_M1_CDNS_7656633918023 $T=59200 80850 0 0 $X=59070 $Y=80770
X546 125 M2_M1_CDNS_7656633918023 $T=59410 91250 0 0 $X=59280 $Y=91170
X547 124 M2_M1_CDNS_7656633918023 $T=61910 97030 0 0 $X=61780 $Y=96950
X548 126 M2_M1_CDNS_7656633918025 $T=-260 63930 0 0 $X=-390 $Y=63800
X549 127 M2_M1_CDNS_7656633918025 $T=3160 97850 0 0 $X=3030 $Y=97720
X550 126 M2_M1_CDNS_7656633918025 $T=6890 63930 0 0 $X=6760 $Y=63800
X551 128 M2_M1_CDNS_7656633918025 $T=12890 59630 0 0 $X=12760 $Y=59500
X552 128 M2_M1_CDNS_7656633918025 $T=12890 64360 0 0 $X=12760 $Y=64230
X553 129 M2_M1_CDNS_7656633918025 $T=18230 63930 0 0 $X=18100 $Y=63800
X554 130 M2_M1_CDNS_7656633918025 $T=20570 64300 0 0 $X=20440 $Y=64170
X555 40 M2_M1_CDNS_7656633918025 $T=21290 80000 0 0 $X=21160 $Y=79870
X556 131 M2_M1_CDNS_7656633918025 $T=27340 60270 0 0 $X=27210 $Y=60140
X557 132 M2_M1_CDNS_7656633918025 $T=28230 63930 0 0 $X=28100 $Y=63800
X558 1 M2_M1_CDNS_7656633918025 $T=30220 101440 0 0 $X=30090 $Y=101310
X559 132 M2_M1_CDNS_7656633918025 $T=30840 58920 0 0 $X=30710 $Y=58790
X560 133 M2_M1_CDNS_7656633918025 $T=31460 59570 0 0 $X=31330 $Y=59440
X561 134 M2_M1_CDNS_7656633918025 $T=37230 64630 0 0 $X=37100 $Y=64500
X562 135 M2_M1_CDNS_7656633918025 $T=40910 64630 0 0 $X=40780 $Y=64500
X563 38 M2_M1_CDNS_7656633918025 $T=50120 100740 0 0 $X=49990 $Y=100610
X564 136 M2_M1_CDNS_7656633918025 $T=53980 60150 0 0 $X=53850 $Y=60020
X565 136 M2_M1_CDNS_7656633918025 $T=54640 63920 0 0 $X=54510 $Y=63790
X566 137 M2_M1_CDNS_7656633918025 $T=55250 65450 0 0 $X=55120 $Y=65320
X567 26 M3_M2_CDNS_7656633918026 $T=230 110810 0 0 $X=-20 $Y=110730
X568 3 M3_M2_CDNS_7656633918026 $T=20130 111380 0 0 $X=19880 $Y=111300
X569 39 M3_M2_CDNS_7656633918026 $T=21380 72640 0 0 $X=21130 $Y=72560
X570 28 M3_M2_CDNS_7656633918026 $T=25910 97510 0 0 $X=25660 $Y=97430
X571 132 M3_M2_CDNS_7656633918026 $T=30840 58920 0 0 $X=30590 $Y=58840
X572 138 M3_M2_CDNS_7656633918026 $T=59210 74060 0 0 $X=58960 $Y=73980
X573 139 M3_M2_CDNS_7656633918026 $T=59230 82660 0 0 $X=58980 $Y=82580
X574 140 M3_M2_CDNS_7656633918026 $T=59260 64440 0 0 $X=59010 $Y=64360
X575 82 M3_M2_CDNS_7656633918027 $T=550 64640 0 0 $X=470 $Y=64390
X576 12 M3_M2_CDNS_7656633918027 $T=2770 110920 0 0 $X=2690 $Y=110670
X577 72 M3_M2_CDNS_7656633918027 $T=7560 120840 0 0 $X=7480 $Y=120590
X578 82 M3_M2_CDNS_7656633918027 $T=11890 64220 0 0 $X=11810 $Y=63970
X579 80 M3_M2_CDNS_7656633918027 $T=17660 71070 0 0 $X=17580 $Y=70820
X580 117 M3_M2_CDNS_7656633918027 $T=22820 59760 0 0 $X=22740 $Y=59510
X581 82 M3_M2_CDNS_7656633918027 $T=23230 64170 0 0 $X=23150 $Y=63920
X582 63 M3_M2_CDNS_7656633918027 $T=25170 89190 0 0 $X=25090 $Y=88940
X583 80 M3_M2_CDNS_7656633918027 $T=28770 71070 0 0 $X=28690 $Y=70820
X584 82 M3_M2_CDNS_7656633918027 $T=34450 64130 0 0 $X=34370 $Y=63880
X585 134 M3_M2_CDNS_7656633918027 $T=35130 59760 0 0 $X=35050 $Y=59510
X586 80 M3_M2_CDNS_7656633918027 $T=40330 79760 0 0 $X=40250 $Y=79510
X587 82 M3_M2_CDNS_7656633918027 $T=45910 64110 0 0 $X=45830 $Y=63860
X588 80 M3_M2_CDNS_7656633918027 $T=51490 79650 0 0 $X=51410 $Y=79400
X589 82 M3_M2_CDNS_7656633918027 $T=57250 64080 0 0 $X=57170 $Y=63830
X590 82 M3_M2_CDNS_7656633918027 $T=59270 49170 0 180 $X=59190 $Y=48920
X591 82 M2_M1_CDNS_7656633918028 $T=550 64640 0 0 $X=470 $Y=64390
X592 12 M2_M1_CDNS_7656633918028 $T=2770 110920 0 0 $X=2690 $Y=110670
X593 72 M2_M1_CDNS_7656633918028 $T=7560 120840 0 0 $X=7480 $Y=120590
X594 82 M2_M1_CDNS_7656633918028 $T=11890 64220 0 0 $X=11810 $Y=63970
X595 80 M2_M1_CDNS_7656633918028 $T=17660 71070 0 0 $X=17580 $Y=70820
X596 82 M2_M1_CDNS_7656633918028 $T=23230 64170 0 0 $X=23150 $Y=63920
X597 63 M2_M1_CDNS_7656633918028 $T=25170 89190 0 0 $X=25090 $Y=88940
X598 80 M2_M1_CDNS_7656633918028 $T=28770 71070 0 0 $X=28690 $Y=70820
X599 82 M2_M1_CDNS_7656633918028 $T=34450 64130 0 0 $X=34370 $Y=63880
X600 80 M2_M1_CDNS_7656633918028 $T=40330 79760 0 0 $X=40250 $Y=79510
X601 82 M2_M1_CDNS_7656633918028 $T=45910 64110 0 0 $X=45830 $Y=63860
X602 80 M2_M1_CDNS_7656633918028 $T=51490 79650 0 0 $X=51410 $Y=79400
X603 82 M2_M1_CDNS_7656633918028 $T=57250 64080 0 0 $X=57170 $Y=63830
X604 127 M3_M2_CDNS_7656633918029 $T=3790 97850 0 0 $X=3660 $Y=97720
X605 126 M3_M2_CDNS_7656633918029 $T=4810 63930 0 0 $X=4680 $Y=63800
X606 117 M3_M2_CDNS_7656633918029 $T=22020 62580 0 0 $X=21890 $Y=62450
X607 133 M3_M2_CDNS_7656633918029 $T=31460 59570 0 0 $X=31330 $Y=59440
X608 134 M3_M2_CDNS_7656633918029 $T=37240 63760 0 0 $X=37110 $Y=63630
X609 14 M4_M3_CDNS_7656633918030 $T=6790 89980 0 0 $X=6420 $Y=89850
X610 25 M4_M3_CDNS_7656633918030 $T=9950 90030 0 0 $X=9580 $Y=89900
X611 20 M4_M3_CDNS_7656633918030 $T=37310 88780 0 0 $X=36940 $Y=88650
X612 27 M4_M3_CDNS_7656633918030 $T=49320 97160 0 0 $X=48950 $Y=97030
X613 69 M3_M2_CDNS_7656633918031 $T=8420 80300 0 0 $X=8290 $Y=80170
X614 66 M3_M2_CDNS_7656633918031 $T=9710 73550 0 0 $X=9580 $Y=73420
X615 35 M3_M2_CDNS_7656633918031 $T=20130 103160 0 0 $X=20000 $Y=103030
X616 9 M3_M2_CDNS_7656633918031 $T=54300 101520 0 0 $X=54170 $Y=101390
X617 14 M3_M2_CDNS_7656633918034 $T=18260 81230 0 0 $X=17890 $Y=81150
X618 59 M3_M2_CDNS_7656633918034 $T=51300 101400 0 0 $X=50930 $Y=101320
X619 64 M3_M2_CDNS_7656633918035 $T=4820 42750 0 0 $X=4740 $Y=42500
X620 4 M3_M2_CDNS_7656633918035 $T=22580 119930 0 0 $X=22500 $Y=119680
X621 127 M4_M3_CDNS_7656633918036 $T=-1050 17310 0 0 $X=-1130 $Y=17060
X622 4 M4_M3_CDNS_7656633918036 $T=22580 119930 0 0 $X=22500 $Y=119680
X623 48 M4_M3_CDNS_7656633918036 $T=37450 101760 0 0 $X=37370 $Y=101510
X624 126 M2_M1_CDNS_7656633918037 $T=-260 57410 0 0 $X=-390 $Y=57280
X625 77 M2_M1_CDNS_7656633918037 $T=870 59200 0 0 $X=740 $Y=59070
X626 141 M2_M1_CDNS_7656633918037 $T=3920 58640 0 0 $X=3790 $Y=58510
X627 126 M2_M1_CDNS_7656633918037 $T=4740 58230 0 0 $X=4610 $Y=58100
X628 81 M2_M1_CDNS_7656633918037 $T=5230 120900 0 0 $X=5100 $Y=120770
X629 141 M2_M1_CDNS_7656633918037 $T=8460 64880 0 0 $X=8330 $Y=64750
X630 142 M2_M1_CDNS_7656633918037 $T=12450 59070 0 0 $X=12320 $Y=58940
X631 142 M2_M1_CDNS_7656633918037 $T=12450 64880 0 0 $X=12320 $Y=64750
X632 130 M2_M1_CDNS_7656633918037 $T=17350 59970 0 0 $X=17220 $Y=59840
X633 129 M2_M1_CDNS_7656633918037 $T=18880 60150 0 0 $X=18750 $Y=60020
X634 117 M2_M1_CDNS_7656633918037 $T=22820 59760 0 0 $X=22690 $Y=59630
X635 131 M2_M1_CDNS_7656633918037 $T=30540 64940 0 0 $X=30410 $Y=64810
X636 133 M2_M1_CDNS_7656633918037 $T=31500 64270 0 0 $X=31370 $Y=64140
X637 134 M2_M1_CDNS_7656633918037 $T=35130 59760 0 0 $X=35000 $Y=59630
X638 143 M2_M1_CDNS_7656633918037 $T=39570 59570 0 0 $X=39440 $Y=59440
X639 143 M2_M1_CDNS_7656633918037 $T=39570 64630 0 0 $X=39440 $Y=64500
X640 94 M2_M1_CDNS_7656633918037 $T=43940 59990 0 0 $X=43810 $Y=59860
X641 135 M2_M1_CDNS_7656633918037 $T=45450 59630 0 0 $X=45320 $Y=59500
X642 98 M2_M1_CDNS_7656633918037 $T=49530 60010 0 0 $X=49400 $Y=59880
X643 122 M2_M1_CDNS_7656633918037 $T=58030 60140 0 0 $X=57900 $Y=60010
X644 137 M2_M1_CDNS_7656633918037 $T=60780 52610 0 0 $X=60650 $Y=52480
X645 144 M2_M1_CDNS_7656633918037 $T=61140 51440 0 0 $X=61010 $Y=51310
X646 144 M2_M1_CDNS_7656633918037 $T=61140 65420 0 0 $X=61010 $Y=65290
X647 145 M3_M2_CDNS_7656633918038 $T=-810 43780 0 0 $X=-940 $Y=43650
X648 146 M3_M2_CDNS_7656633918038 $T=-380 43220 0 0 $X=-510 $Y=43090
X649 132 M3_M2_CDNS_7656633918038 $T=31050 62810 0 0 $X=30920 $Y=62680
X650 147 M3_M2_CDNS_7656633918038 $T=31060 42750 0 0 $X=30930 $Y=42620
X651 133 M3_M2_CDNS_7656633918038 $T=31500 63160 0 0 $X=31370 $Y=63030
X652 140 M3_M2_CDNS_7656633918038 $T=31510 37970 0 0 $X=31380 $Y=37840
X653 138 M3_M2_CDNS_7656633918038 $T=40300 37320 0 0 $X=40170 $Y=37190
X654 139 M3_M2_CDNS_7656633918038 $T=45890 36750 0 0 $X=45760 $Y=36620
X655 147 M3_M2_CDNS_7656633918038 $T=55330 42750 0 0 $X=55200 $Y=42620
X656 138 M2_M1_CDNS_7656633918042 $T=59210 74060 0 0 $X=58960 $Y=73980
X657 139 M2_M1_CDNS_7656633918042 $T=59230 82660 0 0 $X=58980 $Y=82580
X658 74 M3_M2_CDNS_7656633918043 $T=13070 42750 0 0 $X=12820 $Y=42620
X659 75 M3_M2_CDNS_7656633918043 $T=18650 42750 0 0 $X=18400 $Y=42620
X660 74 M4_M3_CDNS_7656633918044 $T=13070 42750 0 0 $X=12820 $Y=42670
X661 148 M4_M3_CDNS_7656633918044 $T=61670 21020 0 0 $X=61420 $Y=20940
X662 149 M4_M3_CDNS_7656633918044 $T=62140 17310 0 0 $X=61890 $Y=17230
X663 64 M5_M4_CDNS_7656633918045 $T=4820 42750 0 0 $X=4740 $Y=42500
X664 65 M5_M4_CDNS_7656633918045 $T=60960 21490 0 0 $X=60880 $Y=21240
X665 65 M7_M6_CDNS_7656633918047 $T=22900 44330 0 0 $X=22770 $Y=44200
X666 148 M7_M6_CDNS_7656633918047 $T=27760 44330 0 0 $X=27630 $Y=44200
X667 148 M5_M4_CDNS_7656633918049 $T=61670 21020 0 0 $X=61420 $Y=20940
X668 149 M5_M4_CDNS_7656633918049 $T=62140 17310 0 0 $X=61890 $Y=17230
X669 148 M3_M2_CDNS_7656633918050 $T=61670 21020 0 0 $X=61420 $Y=20940
X670 149 M3_M2_CDNS_7656633918050 $T=62140 17310 0 0 $X=61890 $Y=17230
X671 65 M7_M6_CDNS_7656633918051 $T=60960 43450 0 0 $X=60830 $Y=43320
X672 148 M7_M6_CDNS_7656633918051 $T=61670 43980 0 0 $X=61540 $Y=43850
X673 149 M7_M6_CDNS_7656633918051 $T=62140 44330 0 0 $X=62010 $Y=44200
X674 148 M6_M5_CDNS_7656633918052 $T=61670 21020 0 0 $X=61420 $Y=20890
X675 149 M6_M5_CDNS_7656633918052 $T=62140 17310 0 0 $X=61890 $Y=17180
X676 65 M6_M5_CDNS_7656633918053 $T=60960 21490 0 0 $X=60880 $Y=21240
X677 127 M3_M2_CDNS_7656633918054 $T=-1050 17310 0 0 $X=-1180 $Y=17060
X678 65 M3_M2_CDNS_7656633918054 $T=60960 21490 0 0 $X=60830 $Y=21240
X679 112 82 76 10 47 80 242 241 598 807
+ 808 599 HAdder $T=-310 72840 0 0 $X=490 $Y=63880
X680 51 82 67 38 9 80 244 243 600 809
+ 810 601 HAdder $T=-310 98645 0 0 $X=490 $Y=89685
X681 77 82 127 76 113 80 246 245 602 811
+ 812 603 HAdder $T=-310 105415 0 0 $X=490 $Y=96455
X682 50 82 78 12 22 80 248 247 604 813
+ 814 605 HAdder $T=-310 112345 0 0 $X=490 $Y=103385
X683 114 82 150 81 32 80 250 249 606 815
+ 816 607 HAdder $T=12750 81440 1 180 $X=6160 $Y=72480
X684 54 82 151 72 50 80 252 251 608 817
+ 818 609 HAdder $T=11030 81440 0 0 $X=11830 $Y=72480
X685 115 82 84 83 152 80 254 253 610 819
+ 820 611 HAdder $T=11030 90040 0 0 $X=11830 $Y=81080
X686 34 82 55 11 46 80 256 255 612 821
+ 822 613 HAdder $T=24090 98645 1 180 $X=17500 $Y=89685
X687 122 82 98 153 97 80 258 257 614 823
+ 824 615 HAdder $T=45050 72840 0 0 $X=45850 $Y=63880
X688 137 82 136 154 100 80 260 259 616 825
+ 826 617 HAdder $T=58110 72840 1 180 $X=51520 $Y=63880
X689 109 82 154 104 101 80 262 261 618 827
+ 828 619 HAdder $T=58110 81440 1 180 $X=51520 $Y=72480
X690 140 82 144 155 109 80 264 263 620 829
+ 830 621 HAdder $T=56390 72840 0 0 $X=57190 $Y=63880
X691 138 82 155 156 106 80 266 265 622 831
+ 832 623 HAdder $T=56390 81440 0 0 $X=57190 $Y=72480
X692 139 82 156 157 111 80 268 267 624 833
+ 834 625 HAdder $T=56390 90040 0 0 $X=57190 $Y=81080
X693 125 82 157 158 110 80 270 269 626 835
+ 836 627 HAdder $T=56390 98640 0 0 $X=57190 $Y=89680
X694 126 141 77 159 82 80 142 145 128 130
+ 146 129 117 65 131 148 132 133 134 149
+ 143 94 64 135 98 75 74 136 122 147
+ 137 144 274 282 286 284 281 310 314 312
+ 309 271 288 292 297 280 316 320 325 273
+ 275 278 279 303 305 306 307 308 WallaceFinalAdder $T=0 42440 0 0 $X=0 $Y=42440
X695 82 69 45 79 49 160 80 335 334 333 FAdder $T=-600 81940 1 0 $X=490 $Y=72480
X696 82 42 41 160 13 36 80 338 337 336 FAdder $T=-600 90540 1 0 $X=490 $Y=81080
X697 82 161 21 162 26 78 80 341 340 339 FAdder $T=-600 109815 0 0 $X=490 $Y=110675
X698 82 126 150 141 66 112 80 344 343 342 FAdder $T=13040 73340 0 180 $X=6160 $Y=63880
X699 82 73 15 57 25 163 80 347 346 345 FAdder $T=13040 90540 0 180 $X=6160 $Y=81080
X700 82 71 43 163 30 16 80 350 349 348 FAdder $T=13040 99145 0 180 $X=6160 $Y=89685
X701 82 14 17 164 53 8 80 353 352 351 FAdder $T=13040 102525 1 180 $X=6160 $Y=103385
X702 82 165 1 166 18 164 80 356 355 354 FAdder $T=13040 109815 1 180 $X=6160 $Y=110675
X703 82 128 151 142 44 114 80 359 358 357 FAdder $T=10740 73340 1 0 $X=11830 $Y=63880
X704 82 20 5 152 48 24 80 362 361 360 FAdder $T=10740 99145 1 0 $X=11830 $Y=89685
X705 82 2 33 167 52 7 80 365 364 363 FAdder $T=10740 102525 0 0 $X=11830 $Y=103385
X706 82 168 19 169 29 167 80 368 367 366 FAdder $T=10740 109815 0 0 $X=11830 $Y=110675
X707 82 129 170 130 39 54 80 371 370 369 FAdder $T=24380 73340 0 180 $X=17500 $Y=63880
X708 82 116 171 170 40 14 80 374 373 372 FAdder $T=24380 81940 0 180 $X=17500 $Y=72480
X709 82 86 67 171 2 60 80 377 376 375 FAdder $T=24380 90540 0 180 $X=17500 $Y=81080
X710 82 63 35 172 58 6 80 380 379 378 FAdder $T=24380 102525 1 180 $X=17500 $Y=103385
X711 82 173 3 174 85 172 80 383 382 381 FAdder $T=24380 109815 1 180 $X=17500 $Y=110675
X712 82 132 175 117 4 116 80 386 385 384 FAdder $T=22080 73340 1 0 $X=23170 $Y=63880
X713 82 118 176 175 23 86 80 389 388 387 FAdder $T=22080 81940 1 0 $X=23170 $Y=72480
X714 82 87 177 176 63 51 80 392 391 390 FAdder $T=22080 90540 1 0 $X=23170 $Y=81080
X715 82 89 31 177 27 28 80 395 394 393 FAdder $T=22080 99145 1 0 $X=23170 $Y=89685
X716 82 133 178 131 79 118 80 398 397 396 FAdder $T=35720 73340 0 180 $X=28840 $Y=63880
X717 82 119 179 178 69 87 80 401 400 399 FAdder $T=35720 81940 0 180 $X=28840 $Y=72480
X718 82 120 180 179 42 89 80 404 403 402 FAdder $T=35720 90540 0 180 $X=28840 $Y=81080
X719 82 56 88 180 103 68 80 407 406 405 FAdder $T=35720 99145 0 180 $X=28840 $Y=89685
X720 82 143 181 134 57 119 80 410 409 408 FAdder $T=33420 73340 1 0 $X=34510 $Y=63880
X721 82 121 182 181 73 120 80 413 412 411 FAdder $T=33420 81940 1 0 $X=34510 $Y=72480
X722 82 93 183 182 71 56 80 416 415 414 FAdder $T=33420 90540 1 0 $X=34510 $Y=81080
X723 82 90 70 183 59 62 80 419 418 417 FAdder $T=33420 99145 1 0 $X=34510 $Y=89685
X724 82 135 184 94 84 121 80 422 421 420 FAdder $T=47060 73340 0 180 $X=40180 $Y=63880
X725 82 97 185 184 115 93 80 425 424 423 FAdder $T=47060 81940 0 180 $X=40180 $Y=72480
X726 82 91 186 185 20 90 80 428 427 426 FAdder $T=47060 90540 0 180 $X=40180 $Y=81080
X727 82 92 105 186 95 37 80 431 430 429 FAdder $T=47060 99145 0 180 $X=40180 $Y=89685
X728 82 100 187 153 55 91 80 434 433 432 FAdder $T=44760 81940 1 0 $X=45850 $Y=72480
X729 82 101 188 187 34 92 80 437 436 435 FAdder $T=44760 90540 1 0 $X=45850 $Y=81080
X730 82 102 107 188 96 99 80 440 439 438 FAdder $T=44760 99145 1 0 $X=45850 $Y=89685
X731 82 106 189 104 61 102 80 443 442 441 FAdder $T=58400 90540 0 180 $X=51520 $Y=81080
X732 82 111 108 189 123 124 80 446 445 444 FAdder $T=58400 99140 0 180 $X=51520 $Y=89680
X733 190 191 192 193 194 195 196 197 198 80
+ 82 62 37 99 124 158 199 200 28 68
+ 70 105 107 108 110 201 9 31 88 103
+ 59 95 96 123 202 60 38 27 36 16
+ 24 46 61 203 8 7 6 35 41 43
+ 5 11 204 22 17 33 52 58 13 30
+ 48 205 32 12 53 19 3 45 15 83
+ 206 47 21 1 18 29 85 49 25 113
+ 10 26 WallaceMultiplier $T=67110 70770 1 180 $X=23170 $Y=101330
X734 162 80 82 66 511 Diver $T=4340 118060 1 90 $X=490 $Y=118790
X735 161 80 82 81 512 Diver $T=7320 118060 1 90 $X=3470 $Y=118790
X736 165 80 82 72 513 Diver $T=5120 118010 0 90 $X=6160 $Y=118740
X737 166 80 82 44 514 Diver $T=8100 118050 0 90 $X=9140 $Y=118780
X738 169 80 82 39 515 Diver $T=15680 118090 1 90 $X=11830 $Y=118820
X739 168 80 82 40 516 Diver $T=18660 118080 1 90 $X=14810 $Y=118810
X740 173 80 82 23 517 Diver $T=16460 118040 0 90 $X=17500 $Y=118770
X741 174 80 82 4 518 Diver $T=19440 118020 0 90 $X=20480 $Y=118750
X742 64 207 82 80 208 209 210 127 74 211
+ 212 213 214 159 75 215 216 217 218 219
+ 220 145 147 146 140 221 222 223 224 225
+ 226 65 138 227 228 229 230 148 139 231
+ 232 233 234 235 236 237 238 149 125 239
+ 240 519 524 536 541 540 538 537 535 534
+ 572 571 576 573 543 549 548 555 554 533
+ 532 578 577 584 583 590 589 522 526 525
+ 529 528 531 530 563 562 565 564 567 566
+ 569 568 570 542 523 740 MAC $T=0 40 0 0 $X=0 $Y=40
M0 511 162 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=1270 $Y=119400 $dt=0
M1 66 511 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=1270 $Y=120330 $dt=0
M2 79 333 45 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=73900 $dt=0
M3 69 333 160 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=75240 $dt=0
M4 333 160 69 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=75650 $dt=0
M5 335 45 334 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=76580 $dt=0
M6 45 334 335 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=76990 $dt=0
M7 333 49 45 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=77400 $dt=0
M8 49 45 333 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=77810 $dt=0
M9 160 336 41 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=82500 $dt=0
M10 42 336 36 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=83840 $dt=0
M11 336 36 42 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=84250 $dt=0
M12 338 41 337 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=85180 $dt=0
M13 41 337 338 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=85590 $dt=0
M14 336 13 41 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=86000 $dt=0
M15 13 41 336 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=86410 $dt=0
M16 339 21 26 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=113855 $dt=0
M17 21 26 339 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=114265 $dt=0
M18 341 340 21 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=114675 $dt=0
M19 340 21 341 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=115085 $dt=0
M20 161 78 339 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=116015 $dt=0
M21 78 339 161 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=116425 $dt=0
M22 21 339 162 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1380 $Y=117765 $dt=0
M23 512 161 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=4250 $Y=119400 $dt=0
M24 81 512 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=4250 $Y=120330 $dt=0
M25 513 165 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=7950 $Y=119350 $dt=0
M26 72 513 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=7950 $Y=120280 $dt=0
M27 141 342 150 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=65300 $dt=0
M28 126 342 112 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=66640 $dt=0
M29 342 112 126 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=67050 $dt=0
M30 344 150 343 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=67980 $dt=0
M31 150 343 344 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=68390 $dt=0
M32 342 66 150 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=68800 $dt=0
M33 66 150 342 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=69210 $dt=0
M34 57 345 15 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=82500 $dt=0
M35 73 345 163 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=83840 $dt=0
M36 345 163 73 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=84250 $dt=0
M37 347 15 346 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=85180 $dt=0
M38 15 346 347 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=85590 $dt=0
M39 345 25 15 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=86000 $dt=0
M40 25 15 345 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=86410 $dt=0
M41 163 348 43 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=91105 $dt=0
M42 71 348 16 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=92445 $dt=0
M43 348 16 71 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=92855 $dt=0
M44 350 43 349 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=93785 $dt=0
M45 43 349 350 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=94195 $dt=0
M46 348 30 43 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=94605 $dt=0
M47 30 43 348 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=95015 $dt=0
M48 351 17 53 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=106565 $dt=0
M49 17 53 351 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=106975 $dt=0
M50 353 352 17 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=107385 $dt=0
M51 352 17 353 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=107795 $dt=0
M52 14 8 351 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=108725 $dt=0
M53 8 351 14 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=109135 $dt=0
M54 17 351 164 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=110475 $dt=0
M55 354 1 18 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=113855 $dt=0
M56 1 18 354 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=114265 $dt=0
M57 356 355 1 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=114675 $dt=0
M58 355 1 356 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=115085 $dt=0
M59 165 164 354 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=116015 $dt=0
M60 164 354 165 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=116425 $dt=0
M61 1 354 166 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=10820 $Y=117765 $dt=0
M62 514 166 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=10930 $Y=119390 $dt=0
M63 44 514 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=10930 $Y=120320 $dt=0
M64 515 169 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=12610 $Y=119430 $dt=0
M65 39 515 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=12610 $Y=120360 $dt=0
M66 142 357 151 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=65300 $dt=0
M67 128 357 114 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=66640 $dt=0
M68 357 114 128 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=67050 $dt=0
M69 359 151 358 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=67980 $dt=0
M70 151 358 359 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=68390 $dt=0
M71 357 44 151 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=68800 $dt=0
M72 44 151 357 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=69210 $dt=0
M73 152 360 5 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=91105 $dt=0
M74 20 360 24 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=92445 $dt=0
M75 360 24 20 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=92855 $dt=0
M76 362 5 361 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=93785 $dt=0
M77 5 361 362 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=94195 $dt=0
M78 360 48 5 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=94605 $dt=0
M79 48 5 360 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=95015 $dt=0
M80 363 33 52 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=106565 $dt=0
M81 33 52 363 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=106975 $dt=0
M82 365 364 33 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=107385 $dt=0
M83 364 33 365 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=107795 $dt=0
M84 2 7 363 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=108725 $dt=0
M85 7 363 2 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=109135 $dt=0
M86 33 363 167 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=110475 $dt=0
M87 366 19 29 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=113855 $dt=0
M88 19 29 366 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=114265 $dt=0
M89 368 367 19 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=114675 $dt=0
M90 367 19 368 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=115085 $dt=0
M91 168 167 366 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=116015 $dt=0
M92 167 366 168 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=116425 $dt=0
M93 19 366 169 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=12720 $Y=117765 $dt=0
M94 516 168 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=15590 $Y=119420 $dt=0
M95 40 516 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=15590 $Y=120350 $dt=0
M96 517 173 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=19290 $Y=119380 $dt=0
M97 23 517 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.682 scb=0.0101159 scc=0.000211679 $X=19290 $Y=120310 $dt=0
M98 130 369 170 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.10357 scb=0.000255666 scc=3.44804e-08 $X=22160 $Y=65300 $dt=0
M99 129 369 54 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=66640 $dt=0
M100 369 54 129 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=67050 $dt=0
M101 371 170 370 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=67980 $dt=0
M102 170 370 371 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=68390 $dt=0
M103 369 39 170 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=68800 $dt=0
M104 39 170 369 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=69210 $dt=0
M105 170 372 171 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=73900 $dt=0
M106 116 372 14 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=75240 $dt=0
M107 372 14 116 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=75650 $dt=0
M108 374 171 373 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=76580 $dt=0
M109 171 373 374 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=76990 $dt=0
M110 372 40 171 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=77400 $dt=0
M111 40 171 372 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=77810 $dt=0
M112 171 375 67 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=82500 $dt=0
M113 86 375 60 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=83840 $dt=0
M114 375 60 86 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=84250 $dt=0
M115 377 67 376 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=85180 $dt=0
M116 67 376 377 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=85590 $dt=0
M117 375 2 67 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=86000 $dt=0
M118 2 67 375 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=86410 $dt=0
M119 378 35 58 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=106565 $dt=0
M120 35 58 378 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=106975 $dt=0
M121 380 379 35 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=107385 $dt=0
M122 379 35 380 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=107795 $dt=0
M123 63 6 378 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=108725 $dt=0
M124 6 378 63 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=109135 $dt=0
M125 35 378 172 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=110475 $dt=0
M126 381 3 85 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=113855 $dt=0
M127 3 85 381 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=114265 $dt=0
M128 383 382 3 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=114675 $dt=0
M129 382 3 383 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=4.11282 scb=0.000306462 scc=1.0989e-07 $X=22160 $Y=115085 $dt=0
M130 173 172 381 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=116015 $dt=0
M131 172 381 173 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=4.52605 scb=0.000482855 scc=2.15388e-07 $X=22160 $Y=116425 $dt=0
M132 3 381 174 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=22160 $Y=117765 $dt=0
M133 518 174 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=22270 $Y=119360 $dt=0
M134 4 518 82 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8263 scb=0.00911451 scc=0.000207374 $X=22270 $Y=120290 $dt=0
M135 117 384 175 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=65300 $dt=0
M136 132 384 116 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=66640 $dt=0
M137 384 116 132 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=67050 $dt=0
M138 386 175 385 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=67980 $dt=0
M139 175 385 386 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=68390 $dt=0
M140 384 4 175 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=68800 $dt=0
M141 4 175 384 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=69210 $dt=0
M142 175 387 176 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=73900 $dt=0
M143 118 387 86 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=75240 $dt=0
M144 387 86 118 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=75650 $dt=0
M145 389 176 388 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=76580 $dt=0
M146 176 388 389 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=76990 $dt=0
M147 387 23 176 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=77400 $dt=0
M148 23 176 387 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=77810 $dt=0
M149 176 390 177 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=82500 $dt=0
M150 87 390 51 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=83840 $dt=0
M151 390 51 87 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=84250 $dt=0
M152 392 177 391 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=85180 $dt=0
M153 177 391 392 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=85590 $dt=0
M154 390 63 177 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=86000 $dt=0
M155 63 177 390 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=86410 $dt=0
M156 177 393 31 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=91105 $dt=0
M157 89 393 28 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=92445 $dt=0
M158 393 28 89 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=92855 $dt=0
M159 395 31 394 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=93785 $dt=0
M160 31 394 395 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=94195 $dt=0
M161 393 27 31 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=94605 $dt=0
M162 27 31 393 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=24060 $Y=95015 $dt=0
M163 131 396 178 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=4.10624 scb=0.000256891 scc=3.49982e-08 $X=33500 $Y=65300 $dt=0
M164 133 396 118 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=66640 $dt=0
M165 396 118 133 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=67050 $dt=0
M166 398 178 397 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=67980 $dt=0
M167 178 397 398 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=68390 $dt=0
M168 396 79 178 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=68800 $dt=0
M169 79 178 396 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=69210 $dt=0
M170 178 399 179 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=73900 $dt=0
M171 119 399 87 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=75240 $dt=0
M172 399 87 119 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=75650 $dt=0
M173 401 179 400 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=76580 $dt=0
M174 179 400 401 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=76990 $dt=0
M175 399 69 179 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=77400 $dt=0
M176 69 179 399 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=77810 $dt=0
M177 179 402 180 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=82500 $dt=0
M178 120 402 89 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=83840 $dt=0
M179 402 89 120 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=84250 $dt=0
M180 404 180 403 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=85180 $dt=0
M181 180 403 404 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=85590 $dt=0
M182 402 42 180 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=86000 $dt=0
M183 42 180 402 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=86410 $dt=0
M184 180 405 88 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=91105 $dt=0
M185 56 405 68 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=92445 $dt=0
M186 405 68 56 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=92855 $dt=0
M187 407 88 406 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=93785 $dt=0
M188 88 406 407 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=94195 $dt=0
M189 405 103 88 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=94605 $dt=0
M190 103 88 405 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=33500 $Y=95015 $dt=0
M191 134 408 181 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.71642 scb=0.000135303 scc=5.64513e-09 $X=35400 $Y=65300 $dt=0
M192 143 408 119 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=66640 $dt=0
M193 408 119 143 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=67050 $dt=0
M194 410 181 409 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=67980 $dt=0
M195 181 409 410 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=68390 $dt=0
M196 408 57 181 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=68800 $dt=0
M197 57 181 408 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=69210 $dt=0
M198 181 411 182 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=73900 $dt=0
M199 121 411 120 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=75240 $dt=0
M200 411 120 121 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=75650 $dt=0
M201 413 182 412 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=76580 $dt=0
M202 182 412 413 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=76990 $dt=0
M203 411 73 182 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=77400 $dt=0
M204 73 182 411 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=77810 $dt=0
M205 182 414 183 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=82500 $dt=0
M206 93 414 56 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=83840 $dt=0
M207 414 56 93 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=84250 $dt=0
M208 416 183 415 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=85180 $dt=0
M209 183 415 416 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=85590 $dt=0
M210 414 71 183 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=86000 $dt=0
M211 71 183 414 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=86410 $dt=0
M212 183 417 70 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=91105 $dt=0
M213 90 417 62 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=92445 $dt=0
M214 417 62 90 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=92855 $dt=0
M215 419 70 418 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=93785 $dt=0
M216 70 418 419 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=94195 $dt=0
M217 417 59 70 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=94605 $dt=0
M218 59 70 417 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=35400 $Y=95015 $dt=0
M219 94 420 184 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=65300 $dt=0
M220 135 420 121 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=66640 $dt=0
M221 420 121 135 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=67050 $dt=0
M222 422 184 421 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=67980 $dt=0
M223 184 421 422 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=68390 $dt=0
M224 420 84 184 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=68800 $dt=0
M225 84 184 420 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=69210 $dt=0
M226 184 423 185 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=73900 $dt=0
M227 97 423 93 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=75240 $dt=0
M228 423 93 97 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=75650 $dt=0
M229 425 185 424 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=76580 $dt=0
M230 185 424 425 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=76990 $dt=0
M231 423 115 185 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=77400 $dt=0
M232 115 185 423 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=77810 $dt=0
M233 185 426 186 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=82500 $dt=0
M234 91 426 90 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=83840 $dt=0
M235 426 90 91 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=84250 $dt=0
M236 428 186 427 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=85180 $dt=0
M237 186 427 428 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=85590 $dt=0
M238 426 20 186 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=86000 $dt=0
M239 20 186 426 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=86410 $dt=0
M240 186 429 105 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=91105 $dt=0
M241 92 429 37 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=92445 $dt=0
M242 429 37 92 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=92855 $dt=0
M243 431 105 430 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=93785 $dt=0
M244 105 430 431 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=94195 $dt=0
M245 429 95 105 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=94605 $dt=0
M246 95 105 429 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=44840 $Y=95015 $dt=0
M247 153 432 187 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=73900 $dt=0
M248 100 432 91 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=75240 $dt=0
M249 432 91 100 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=75650 $dt=0
M250 434 187 433 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=76580 $dt=0
M251 187 433 434 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=76990 $dt=0
M252 432 55 187 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=77400 $dt=0
M253 55 187 432 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=77810 $dt=0
M254 187 435 188 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=82500 $dt=0
M255 101 435 92 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=83840 $dt=0
M256 435 92 101 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=84250 $dt=0
M257 437 188 436 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=85180 $dt=0
M258 188 436 437 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=85590 $dt=0
M259 435 34 188 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=86000 $dt=0
M260 34 188 435 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=86410 $dt=0
M261 188 438 107 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=91105 $dt=0
M262 102 438 99 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=92445 $dt=0
M263 438 99 102 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=92855 $dt=0
M264 440 107 439 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=93785 $dt=0
M265 107 439 440 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=94195 $dt=0
M266 438 96 107 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=94605 $dt=0
M267 96 107 438 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=46740 $Y=95015 $dt=0
M268 104 441 189 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=82500 $dt=0
M269 106 441 102 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=83840 $dt=0
M270 441 102 106 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=84250 $dt=0
M271 443 189 442 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=85180 $dt=0
M272 189 442 443 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=85590 $dt=0
M273 441 61 189 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=86000 $dt=0
M274 61 189 441 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=86410 $dt=0
M275 189 444 108 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=91100 $dt=0
M276 111 444 124 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=92440 $dt=0
M277 444 124 111 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=92850 $dt=0
M278 446 108 445 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=93780 $dt=0
M279 108 445 446 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=94190 $dt=0
M280 444 123 108 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=94600 $dt=0
M281 123 108 444 82 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=56180 $Y=95010 $dt=0
M282 511 162 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=2280 $Y=119400 $dt=1
M283 66 511 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=2280 $Y=120330 $dt=1
M284 79 333 160 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=4830 $Y=73900 $dt=1
M285 160 336 36 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=4830 $Y=82500 $dt=1
M286 78 339 162 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=4830 $Y=117765 $dt=1
M287 808 242 76 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=65950 $dt=1
M288 80 241 808 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=5210 $Y=66160 $dt=1
M289 80 241 807 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=5210 $Y=67090 $dt=1
M290 807 242 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=5210 $Y=67500 $dt=1
M291 112 47 807 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=67910 $dt=1
M292 807 10 112 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=68320 $dt=1
M293 80 10 241 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5210 $Y=69250 $dt=1
M294 80 47 242 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=70180 $dt=1
M295 810 244 67 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=91755 $dt=1
M296 80 243 810 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=5210 $Y=91965 $dt=1
M297 80 243 809 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=5210 $Y=92895 $dt=1
M298 809 244 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=5210 $Y=93305 $dt=1
M299 51 9 809 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=93715 $dt=1
M300 809 38 51 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=94125 $dt=1
M301 80 38 243 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5210 $Y=95055 $dt=1
M302 80 9 244 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=95985 $dt=1
M303 812 246 127 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5210 $Y=98525 $dt=1
M304 80 245 812 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=5210 $Y=98735 $dt=1
M305 80 245 811 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=5210 $Y=99665 $dt=1
M306 811 246 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=5210 $Y=100075 $dt=1
M307 77 113 811 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=5210 $Y=100485 $dt=1
M308 811 76 77 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=5210 $Y=100895 $dt=1
M309 80 76 245 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=5210 $Y=101825 $dt=1
M310 80 113 246 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5210 $Y=102755 $dt=1
M311 814 248 78 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=105455 $dt=1
M312 80 247 814 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=5210 $Y=105665 $dt=1
M313 80 247 813 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=5210 $Y=106595 $dt=1
M314 813 248 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=5210 $Y=107005 $dt=1
M315 50 22 813 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=107415 $dt=1
M316 813 12 50 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5210 $Y=107825 $dt=1
M317 80 12 247 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=5210 $Y=108755 $dt=1
M318 80 22 248 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=5210 $Y=109685 $dt=1
M319 512 161 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=5260 $Y=119400 $dt=1
M320 81 512 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=5260 $Y=120330 $dt=1
M321 513 165 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=6940 $Y=119350 $dt=1
M322 72 513 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=6940 $Y=120280 $dt=1
M323 816 250 150 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=6990 $Y=74550 $dt=1
M324 80 249 816 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=6990 $Y=74760 $dt=1
M325 80 249 815 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=6990 $Y=75690 $dt=1
M326 815 250 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=6990 $Y=76100 $dt=1
M327 114 32 815 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6990 $Y=76510 $dt=1
M328 815 81 114 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6990 $Y=76920 $dt=1
M329 80 81 249 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=6990 $Y=77850 $dt=1
M330 80 32 250 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=6990 $Y=78780 $dt=1
M331 141 342 112 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=7370 $Y=65300 $dt=1
M332 57 345 163 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=7370 $Y=82500 $dt=1
M333 163 348 16 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=7370 $Y=91105 $dt=1
M334 8 351 164 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=7370 $Y=110475 $dt=1
M335 164 354 166 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=7370 $Y=117765 $dt=1
M336 514 166 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=9920 $Y=119390 $dt=1
M337 44 514 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=9920 $Y=120320 $dt=1
M338 515 169 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=13620 $Y=119430 $dt=1
M339 39 515 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=13620 $Y=120360 $dt=1
M340 142 357 114 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=16170 $Y=65300 $dt=1
M341 152 360 24 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=16170 $Y=91105 $dt=1
M342 7 363 167 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=16170 $Y=110475 $dt=1
M343 167 366 169 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=16170 $Y=117765 $dt=1
M344 818 252 151 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=74550 $dt=1
M345 80 251 818 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=16550 $Y=74760 $dt=1
M346 80 251 817 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=16550 $Y=75690 $dt=1
M347 817 252 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=16550 $Y=76100 $dt=1
M348 54 50 817 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=76510 $dt=1
M349 817 72 54 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=76920 $dt=1
M350 80 72 251 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=16550 $Y=77850 $dt=1
M351 80 50 252 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=78780 $dt=1
M352 820 254 84 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=83150 $dt=1
M353 80 253 820 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=16550 $Y=83360 $dt=1
M354 80 253 819 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=16550 $Y=84290 $dt=1
M355 819 254 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=16550 $Y=84700 $dt=1
M356 115 152 819 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=85110 $dt=1
M357 819 83 115 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16550 $Y=85520 $dt=1
M358 80 83 253 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=16550 $Y=86450 $dt=1
M359 80 152 254 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=16550 $Y=87380 $dt=1
M360 516 168 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=16600 $Y=119420 $dt=1
M361 40 516 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=16600 $Y=120350 $dt=1
M362 517 173 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=18280 $Y=119380 $dt=1
M363 23 517 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=116.208 scb=0.059453 scc=0.0138338 $X=18280 $Y=120310 $dt=1
M364 822 256 55 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=18330 $Y=91755 $dt=1
M365 80 255 822 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=18330 $Y=91965 $dt=1
M366 80 255 821 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=18330 $Y=92895 $dt=1
M367 821 256 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=18330 $Y=93305 $dt=1
M368 34 46 821 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=18330 $Y=93715 $dt=1
M369 821 11 34 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=18330 $Y=94125 $dt=1
M370 80 11 255 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=18330 $Y=95055 $dt=1
M371 80 46 256 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=18330 $Y=95985 $dt=1
M372 130 369 54 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=18710 $Y=65300 $dt=1
M373 170 372 14 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=18710 $Y=73900 $dt=1
M374 171 375 60 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=18710 $Y=82500 $dt=1
M375 6 378 172 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=18710 $Y=110475 $dt=1
M376 172 381 174 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=18710 $Y=117765 $dt=1
M377 518 174 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=21260 $Y=119360 $dt=1
M378 4 518 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=121.853 scb=0.0675097 scc=0.0140235 $X=21260 $Y=120290 $dt=1
M379 117 384 116 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=65300 $dt=1
M380 175 387 86 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=73900 $dt=1
M381 176 390 51 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=82500 $dt=1
M382 177 393 28 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=27510 $Y=91105 $dt=1
M383 131 396 118 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=65300 $dt=1
M384 178 399 87 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=73900 $dt=1
M385 179 402 89 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=82500 $dt=1
M386 180 405 68 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=30050 $Y=91105 $dt=1
M387 134 408 119 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=65300 $dt=1
M388 181 411 120 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=73900 $dt=1
M389 182 414 56 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=82500 $dt=1
M390 183 417 62 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=38850 $Y=91105 $dt=1
M391 94 420 121 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=65300 $dt=1
M392 184 423 93 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=73900 $dt=1
M393 185 426 90 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=82500 $dt=1
M394 186 429 37 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=41390 $Y=91105 $dt=1
M395 153 432 91 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=114.504 scb=0.0583006 scc=0.0134535 $X=50190 $Y=73900 $dt=1
M396 187 435 92 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=50190 $Y=82500 $dt=1
M397 188 438 99 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=50190 $Y=91105 $dt=1
M398 824 258 98 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=50570 $Y=65950 $dt=1
M399 80 257 824 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.901 scb=0.0471116 scc=0.0116656 $X=50570 $Y=66160 $dt=1
M400 80 257 823 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.1268 scb=0.0349743 scc=0.0111863 $X=50570 $Y=67090 $dt=1
M401 823 258 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.5388 scb=0.0347327 scc=0.0111862 $X=50570 $Y=67500 $dt=1
M402 122 97 823 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=50570 $Y=67910 $dt=1
M403 823 153 122 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=50570 $Y=68320 $dt=1
M404 80 153 257 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.6513 scb=0.0354006 scc=0.011187 $X=50570 $Y=69250 $dt=1
M405 80 97 258 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=50570 $Y=70180 $dt=1
M406 826 260 136 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=52350 $Y=65950 $dt=1
M407 80 259 826 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.901 scb=0.0471116 scc=0.0116656 $X=52350 $Y=66160 $dt=1
M408 80 259 825 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.1268 scb=0.0349743 scc=0.0111863 $X=52350 $Y=67090 $dt=1
M409 825 260 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.5388 scb=0.0347327 scc=0.0111862 $X=52350 $Y=67500 $dt=1
M410 137 100 825 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=52350 $Y=67910 $dt=1
M411 825 154 137 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.4902 scb=0.0347233 scc=0.0111862 $X=52350 $Y=68320 $dt=1
M412 80 154 259 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.6513 scb=0.0354006 scc=0.011187 $X=52350 $Y=69250 $dt=1
M413 80 100 260 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.941 scb=0.0587511 scc=0.0138331 $X=52350 $Y=70180 $dt=1
M414 828 262 154 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52350 $Y=74550 $dt=1
M415 80 261 828 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=52350 $Y=74760 $dt=1
M416 80 261 827 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=52350 $Y=75690 $dt=1
M417 827 262 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=95.4479 scb=0.0347169 scc=0.0111862 $X=52350 $Y=76100 $dt=1
M418 109 101 827 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52350 $Y=76510 $dt=1
M419 827 104 109 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=52350 $Y=76920 $dt=1
M420 80 104 261 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.5604 scb=0.0353848 scc=0.011187 $X=52350 $Y=77850 $dt=1
M421 80 101 262 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=114.851 scb=0.0587353 scc=0.0138331 $X=52350 $Y=78780 $dt=1
M422 104 441 102 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52730 $Y=82500 $dt=1
M423 189 444 124 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=113.117 scb=0.0574313 scc=0.0134521 $X=52730 $Y=91100 $dt=1
M424 830 264 144 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=65950 $dt=1
M425 80 263 830 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=66160 $dt=1
M426 80 263 829 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=67090 $dt=1
M427 829 264 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=67500 $dt=1
M428 140 109 829 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=67910 $dt=1
M429 829 155 140 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=68320 $dt=1
M430 80 155 263 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=69250 $dt=1
M431 80 109 264 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=70180 $dt=1
M432 832 266 155 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=74550 $dt=1
M433 80 265 832 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=74760 $dt=1
M434 80 265 831 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=75690 $dt=1
M435 831 266 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=76100 $dt=1
M436 138 106 831 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=76510 $dt=1
M437 831 156 138 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=76920 $dt=1
M438 80 156 265 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=77850 $dt=1
M439 80 106 266 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=78780 $dt=1
M440 834 268 156 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=83150 $dt=1
M441 80 267 834 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=83360 $dt=1
M442 80 267 833 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=84290 $dt=1
M443 833 268 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=84700 $dt=1
M444 139 111 833 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=85110 $dt=1
M445 833 157 139 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=85520 $dt=1
M446 80 157 267 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=86450 $dt=1
M447 80 111 268 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=87380 $dt=1
M448 836 270 157 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=91750 $dt=1
M449 80 269 836 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=107.421 scb=0.0513211 scc=0.0117083 $X=61910 $Y=91960 $dt=1
M450 80 269 835 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=99.647 scb=0.0391838 scc=0.011229 $X=61910 $Y=92890 $dt=1
M451 835 270 80 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=99.0591 scb=0.0389422 scc=0.0112289 $X=61910 $Y=93300 $dt=1
M452 125 110 835 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=93710 $dt=1
M453 835 158 125 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=99.0105 scb=0.0389328 scc=0.0112289 $X=61910 $Y=94120 $dt=1
M454 80 158 269 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=61910 $Y=95050 $dt=1
M455 80 110 270 80 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=61910 $Y=95980 $dt=1
.ends WallaceProjectMAC
