* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : WallaceFinalAdder                            *
* Netlisted  : Thu Dec 11 09:02:36 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750680                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750680 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750680

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750681                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750681 1 2 3
** N=4 EP=3 FDC=1
M0 2 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765461750681

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750682                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750682 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750682

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750685                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750685 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750685

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND b a Vdd gnd Vout 6
*.DEVICECLIMB
** N=7 EP=6 FDC=4
X7 gnd Vout 6 nmos1v_CDNS_765461750680 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X8 Vdd Vout 6 pmos1v_CDNS_765461750681 $T=4560 -1510 0 0 $X=3880 $Y=-1710
X9 gnd b 7 nmos1v_CDNS_765461750682 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X12 6 a 7 gnd nmos1v_CDNS_765461750685 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750687                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750687 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750687

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR a vdd gnd f b 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X20 gnd gnd a 6 nmos1v_CDNS_765461750687 $T=420 800 0 0 $X=0 $Y=240
X21 f gnd b 6 nmos1v_CDNS_765461750687 $T=1440 800 1 180 $X=930 $Y=240
X22 f gnd 7 a nmos1v_CDNS_765461750687 $T=2280 800 0 0 $X=1860 $Y=240
X23 gnd gnd b 7 nmos1v_CDNS_765461750687 $T=3300 800 1 180 $X=2790 $Y=240
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765461750688                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765461750688 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765461750688

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765461750689                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765461750689 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765461750689

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506810                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506810 1 2 3
** N=4 EP=3 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506810

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506811                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506811 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506811

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506812                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506812 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506812

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506814                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506814 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506814

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506815                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506815 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506815

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506816                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506816 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506816

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506817                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506817 1 2 3
** N=4 EP=3 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506817

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506818                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506818 1 2 3 5
** N=5 EP=4 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506818

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder sum gnd carry a b vdd
** N=12 EP=6 FDC=16
X19 gnd gnd a 8 nmos1v_CDNS_765461750687 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X20 gnd gnd b 7 nmos1v_CDNS_765461750687 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X36 sum b 9 vdd pmos1v_CDNS_765461750688 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 gnd 7 carry nmos1v_CDNS_765461750689 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 9 vdd 7 pmos1v_CDNS_7654617506810 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 vdd 8 11 pmos1v_CDNS_7654617506811 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 carry 7 11 vdd pmos1v_CDNS_7654617506812 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X43 10 7 gnd nmos1v_CDNS_7654617506814 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 a sum 12 gnd nmos1v_CDNS_7654617506815 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 gnd b 12 nmos1v_CDNS_7654617506816 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 9 8 vdd pmos1v_CDNS_7654617506817 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 9 a sum vdd pmos1v_CDNS_7654617506818 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 gnd 8 carry gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 10 8 sum gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M2 vdd a 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=5520 $Y=-3590 $dt=1
M3 vdd b 7 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5520 $Y=-2660 $dt=1
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7654617506819                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7654617506819 1 2 3 4
** N=5 EP=4 FDC=1
M0 4 3 1 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7654617506819

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7654617506820                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7654617506820 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7654617506820

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic p1 g1 c0 vdd gnd p2 g2 cout1 p3 g3
+ cout2 p4 cout3 g4 cout4 19 29
*.DEVICECLIMB
** N=39 EP=17 FDC=54
X91 gnd gnd p1 30 nmos1v_CDNS_765461750687 $T=1030 800 0 0 $X=610 $Y=240
X92 30 gnd c0 16 nmos1v_CDNS_765461750687 $T=1960 800 0 0 $X=1540 $Y=240
X93 gnd gnd p2 31 nmos1v_CDNS_765461750687 $T=4750 800 0 0 $X=4330 $Y=240
X94 31 gnd g1 17 nmos1v_CDNS_765461750687 $T=7540 800 0 0 $X=7120 $Y=240
X95 gnd gnd g2 17 nmos1v_CDNS_765461750687 $T=8560 800 1 180 $X=8050 $Y=240
X96 gnd gnd 17 cout2 nmos1v_CDNS_765461750687 $T=9400 800 0 0 $X=8980 $Y=240
X97 32 gnd p1 33 nmos1v_CDNS_765461750687 $T=12190 800 0 0 $X=11770 $Y=240
X98 33 gnd c0 18 nmos1v_CDNS_765461750687 $T=13120 800 0 0 $X=12700 $Y=240
X99 34 gnd g2 18 nmos1v_CDNS_765461750687 $T=14980 800 0 0 $X=14560 $Y=240
X100 gnd gnd g3 18 nmos1v_CDNS_765461750687 $T=16000 800 1 180 $X=15490 $Y=240
X101 gnd gnd 18 cout3 nmos1v_CDNS_765461750687 $T=16840 800 0 0 $X=16420 $Y=240
X102 35 gnd p3 36 nmos1v_CDNS_765461750687 $T=18700 800 0 0 $X=18280 $Y=240
X103 36 gnd g2 19 nmos1v_CDNS_765461750687 $T=23350 800 0 0 $X=22930 $Y=240
X104 gnd gnd 19 cout4 nmos1v_CDNS_765461750687 $T=26140 800 0 0 $X=25720 $Y=240
X326 vdd vdd p1 16 pmos1v_CDNS_7654617506819 $T=1030 8610 1 0 $X=610 $Y=8170
X327 20 vdd c0 16 pmos1v_CDNS_7654617506819 $T=2050 8610 0 180 $X=1540 $Y=8170
X328 22 vdd p1 17 pmos1v_CDNS_7654617506819 $T=5770 8610 0 180 $X=5260 $Y=8170
X329 vdd vdd 18 cout3 pmos1v_CDNS_7654617506819 $T=16840 8610 1 0 $X=16420 $Y=8170
X330 29 vdd p3 19 pmos1v_CDNS_7654617506819 $T=18790 8610 0 180 $X=18280 $Y=8170
X331 28 vdd c0 19 pmos1v_CDNS_7654617506819 $T=21580 8610 0 180 $X=21070 $Y=8170
X332 29 vdd g3 26 pmos1v_CDNS_7654617506819 $T=24370 8610 0 180 $X=23860 $Y=8170
X333 gnd gnd g1 16 nmos1v_CDNS_7654617506820 $T=2980 1040 0 180 $X=2470 $Y=240
X334 gnd gnd 16 cout1 nmos1v_CDNS_7654617506820 $T=3820 1040 1 0 $X=3400 $Y=240
X335 31 gnd p1 37 nmos1v_CDNS_7654617506820 $T=5680 1040 1 0 $X=5260 $Y=240
X336 37 gnd c0 17 nmos1v_CDNS_7654617506820 $T=6610 1040 1 0 $X=6190 $Y=240
X337 gnd gnd p3 34 nmos1v_CDNS_7654617506820 $T=10330 1040 1 0 $X=9910 $Y=240
X338 34 gnd p2 32 nmos1v_CDNS_7654617506820 $T=11260 1040 1 0 $X=10840 $Y=240
X339 32 gnd g1 18 nmos1v_CDNS_7654617506820 $T=14050 1040 1 0 $X=13630 $Y=240
X340 gnd gnd p4 35 nmos1v_CDNS_7654617506820 $T=17770 1040 1 0 $X=17350 $Y=240
X341 36 gnd p2 38 nmos1v_CDNS_7654617506820 $T=19630 1040 1 0 $X=19210 $Y=240
X342 38 gnd p1 39 nmos1v_CDNS_7654617506820 $T=20560 1040 1 0 $X=20140 $Y=240
X343 39 gnd c0 19 nmos1v_CDNS_7654617506820 $T=21490 1040 1 0 $X=21070 $Y=240
X344 38 gnd g1 19 nmos1v_CDNS_7654617506820 $T=22420 1040 1 0 $X=22000 $Y=240
X345 35 gnd g3 19 nmos1v_CDNS_7654617506820 $T=24280 1040 1 0 $X=23860 $Y=240
X346 gnd gnd g4 19 nmos1v_CDNS_7654617506820 $T=25300 1040 0 180 $X=24790 $Y=240
M0 vdd g1 20 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M1 cout1 16 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M2 17 p2 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M3 21 c0 17 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M4 22 g1 21 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M5 vdd g2 22 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M6 cout2 17 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M7 18 p3 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M8 23 p2 18 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M9 24 p1 18 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M10 25 c0 18 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M11 24 g1 25 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M12 23 g2 24 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M13 vdd g3 23 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M14 19 p4 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M15 26 p2 19 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M16 27 p1 19 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M17 27 g1 28 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M18 26 g2 27 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: WallaceFinalAdder                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt WallaceFinalAdder aout<10> aout<11> aout<12> aout<13> aout<14> aout<5> aout<6> aout<7> aout<8> aout<9>
+ bout<10> bout<11> bout<12> bout<13> bout<14> bout<5> bout<6> bout<7> bout<8> bout<9>
+ gnd s<10> s<11> s<12> s<13> s<14> s<5> s<6> s<7> s<8>
+ s<9> vdd
** N=164 EP=32 FDC=320
X100 bout<13> aout<13> vdd gnd 18 59 AND $T=3670 21910 0 0 $X=4740 $Y=18810
X101 bout<12> aout<12> vdd gnd 19 60 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X102 bout<11> aout<11> vdd gnd 20 61 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X103 bout<10> aout<10> vdd gnd 21 62 AND $T=32210 21910 1 180 $X=26960 $Y=18810
X104 bout<9> aout<9> vdd gnd 22 63 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X105 bout<8> aout<8> vdd gnd 23 64 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X106 bout<7> aout<7> vdd gnd 24 65 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X107 bout<6> aout<6> vdd gnd 25 66 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X108 aout<14> vdd gnd 1 bout<14> 103 67 XOR $T=530 18810 1 0 $X=530 $Y=14110
X109 26 vdd gnd s<14> 1 104 68 XOR $T=640 4700 1 0 $X=640 $Y=0
X110 aout<13> vdd gnd 2 bout<13> 105 69 XOR $T=4740 18810 1 0 $X=4740 $Y=14110
X111 27 vdd gnd s<13> 2 106 70 XOR $T=9740 4700 0 180 $X=6020 $Y=0
X112 28 vdd gnd s<12> 3 107 71 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X113 aout<12> vdd gnd 3 bout<12> 108 72 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X114 29 vdd gnd s<11> 4 109 73 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X115 aout<11> vdd gnd 4 bout<11> 110 74 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X116 30 vdd gnd s<10> 5 111 75 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X117 aout<10> vdd gnd 5 bout<10> 112 76 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X118 aout<9> vdd gnd 6 bout<9> 113 77 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X119 31 vdd gnd s<9> 6 114 78 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X120 32 vdd gnd s<8> 7 115 79 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X121 aout<8> vdd gnd 7 bout<8> 116 80 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X122 33 vdd gnd s<7> 8 117 81 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X123 aout<7> vdd gnd 8 bout<7> 118 82 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X124 54 vdd gnd s<6> 9 119 83 XOR $T=49650 4700 1 0 $X=49650 $Y=0
X125 aout<6> vdd gnd 9 bout<6> 120 84 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X126 s<5> gnd 54 aout<5> bout<5> vdd HAdder $T=62720 6180 1 90 $X=53760 $Y=6980
X127 5 21 30 vdd gnd 4 20 29 3 19
+ 28 2 27 18 26 90 151 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X128 9 25 54 vdd gnd 8 24 33 7 23
+ 32 6 31 22 30 94 161 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
M0 vdd 90 26 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M1 103 aout<14> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=103.81 scb=0.0470958 scc=0.0116656 $X=950 $Y=14910 $dt=1
M2 104 26 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=800 $dt=1
M3 151 18 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M4 1 bout<14> aout<14> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.0359 scb=0.0349585 scc=0.0111863 $X=1880 $Y=14910 $dt=1
M5 s<14> 1 26 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=800 $dt=1
M6 103 67 1 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=2810 $Y=14910 $dt=1
M7 104 68 s<14> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=800 $dt=1
M8 vdd bout<14> 67 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=3740 $Y=14910 $dt=1
M9 vdd 1 68 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=800 $dt=1
M10 105 aout<13> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=14910 $dt=1
M11 59 aout<13> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=20590 $dt=1
M12 vdd bout<13> 59 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=20590 $dt=1
M13 2 bout<13> aout<13> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=14910 $dt=1
M14 70 2 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=800 $dt=1
M15 105 69 2 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=14910 $dt=1
M16 s<13> 70 106 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=800 $dt=1
M17 vdd bout<13> 69 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=14910 $dt=1
M18 27 2 s<13> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=800 $dt=1
M19 vdd 27 106 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=800 $dt=1
M20 71 3 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M21 108 aout<12> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M22 60 aout<12> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=20590 $dt=1
M23 vdd bout<12> 60 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=20590 $dt=1
M24 s<12> 71 107 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M25 3 bout<12> aout<12> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M26 28 3 s<12> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M27 108 72 3 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M28 vdd 28 107 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M29 vdd bout<12> 72 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M30 73 4 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M31 110 aout<11> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M32 61 aout<11> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=20590 $dt=1
M33 s<11> 73 109 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M34 vdd bout<11> 61 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=20590 $dt=1
M35 4 bout<11> aout<11> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M36 29 4 s<11> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M37 110 74 4 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M38 vdd 29 109 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M39 vdd bout<11> 74 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M40 75 5 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M41 s<10> 75 111 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M42 30 5 s<10> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M43 vdd 30 111 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M44 vdd 94 30 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M45 76 bout<10> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M46 161 22 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M47 5 76 112 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M48 aout<10> bout<10> 5 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M49 62 bout<10> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29780 $Y=20590 $dt=1
M50 vdd aout<10> 62 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30190 $Y=20590 $dt=1
M51 vdd aout<10> 112 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M52 113 aout<9> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M53 63 aout<9> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=20590 $dt=1
M54 vdd bout<9> 63 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=20590 $dt=1
M55 6 bout<9> aout<9> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M56 78 6 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M57 113 77 6 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M58 s<9> 78 114 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M59 vdd bout<9> 77 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M60 31 6 s<9> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M61 vdd 31 114 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M62 79 7 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M63 116 aout<8> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M64 64 aout<8> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=20590 $dt=1
M65 vdd bout<8> 64 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=20590 $dt=1
M66 s<8> 79 115 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M67 7 bout<8> aout<8> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M68 32 7 s<8> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M69 116 80 7 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M70 vdd 32 115 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M71 vdd bout<8> 80 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M72 81 8 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M73 118 aout<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M74 65 aout<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=20590 $dt=1
M75 s<7> 81 117 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M76 vdd bout<7> 65 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=20590 $dt=1
M77 8 bout<7> aout<7> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M78 33 8 s<7> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=48010 $Y=800 $dt=1
M79 118 82 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M80 vdd 33 117 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=48940 $Y=800 $dt=1
M81 vdd bout<7> 82 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M82 119 54 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=50070 $Y=800 $dt=1
M83 s<6> 9 54 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=51000 $Y=800 $dt=1
M84 119 83 s<6> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=51930 $Y=800 $dt=1
M85 vdd 9 83 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=52860 $Y=800 $dt=1
M86 84 bout<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M87 9 84 120 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M88 aout<6> bout<6> 9 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M89 66 bout<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=20590 $dt=1
M90 vdd aout<6> 66 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=20590 $dt=1
M91 vdd aout<6> 120 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
.ends WallaceFinalAdder
