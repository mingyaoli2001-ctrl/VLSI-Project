* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : HAdder                                       *
* Netlisted  : Sat Dec  6 20:20:42 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765070438331                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765070438331 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765070438331

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765070438332                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765070438332 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765070438332

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765070438333                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765070438333 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765070438333

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765070438334                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765070438334 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765070438334

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_765070438335                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_765070438335 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_765070438335

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_765070438336                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_765070438336 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_765070438336

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765070438330                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765070438330 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends pmos1v_CDNS_765070438330

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765070438331                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765070438331 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=100.294 scb=0.0411762 scc=0.0112988 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765070438331

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765070438332                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765070438332 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765070438332

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765070438333                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765070438333 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=100.342 scb=0.0411856 scc=0.0112988 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765070438333

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765070438334                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765070438334 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=108.704 scb=0.0535645 scc=0.0117782 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765070438334

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765070438335                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765070438335 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=119.745 scb=0.065204 scc=0.0139457 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765070438335

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765070438336                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765070438336 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_765070438336

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765070438337                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765070438337 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765070438337

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765070438338                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765070438338 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765070438338

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765070438339                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765070438339 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765070438339

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7650704383310                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7650704383310 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=100.93 scb=0.0414272 scc=0.0112989 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7650704383310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7650704383311                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7650704383311 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=100.294 scb=0.0411762 scc=0.0112988 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7650704383311

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7650704383312                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7650704383312 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7650704383312

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder 3 7 10 9 5 8
** N=12 EP=6 FDC=16
X0 1 M2_M1_CDNS_765070438331 $T=1300 -5710 0 270 $X=1170 $Y=-5840
X1 1 M2_M1_CDNS_765070438331 $T=1300 -4270 0 270 $X=1170 $Y=-4400
X2 2 M2_M1_CDNS_765070438332 $T=2340 -4370 0 90 $X=2090 $Y=-4450
X3 2 M2_M1_CDNS_765070438332 $T=2930 -6480 0 90 $X=2680 $Y=-6560
X4 2 M2_M1_CDNS_765070438332 $T=2950 -5710 0 90 $X=2700 $Y=-5790
X5 3 M2_M1_CDNS_765070438332 $T=3490 -4140 0 90 $X=3240 $Y=-4220
X6 3 M2_M1_CDNS_765070438332 $T=3500 -3460 0 90 $X=3250 $Y=-3540
X7 4 M2_M1_CDNS_765070438332 $T=5640 -5920 0 90 $X=5390 $Y=-6000
X8 4 M2_M1_CDNS_765070438332 $T=5640 -5080 0 90 $X=5390 $Y=-5160
X9 4 M2_M1_CDNS_765070438332 $T=5640 -4300 0 90 $X=5390 $Y=-4380
X10 5 M2_M1_CDNS_765070438333 $T=2220 -7390 0 90 $X=2090 $Y=-7470
X11 5 M2_M1_CDNS_765070438333 $T=2220 -4680 0 90 $X=2090 $Y=-4760
X12 6 M2_M1_CDNS_765070438333 $T=4200 -2840 0 90 $X=4070 $Y=-2920
X13 2 M2_M1_CDNS_765070438333 $T=4570 -3920 0 90 $X=4440 $Y=-4000
X14 2 M1_PO_CDNS_765070438334 $T=2340 -4370 0 90 $X=2090 $Y=-4470
X15 2 M1_PO_CDNS_765070438334 $T=2930 -6480 0 90 $X=2680 $Y=-6580
X16 2 M1_PO_CDNS_765070438334 $T=2950 -5710 0 90 $X=2700 $Y=-5810
X17 3 M1_PO_CDNS_765070438334 $T=3490 -4140 0 90 $X=3240 $Y=-4240
X18 3 M1_PO_CDNS_765070438334 $T=3500 -3460 0 90 $X=3250 $Y=-3560
X19 3 M2_M1_CDNS_765070438335 $T=3500 -4810 0 0 $X=3250 $Y=-4940
X20 3 M2_M1_CDNS_765070438335 $T=3500 -1930 0 0 $X=3250 $Y=-2060
X21 6 M2_M1_CDNS_765070438335 $T=4210 -6730 0 0 $X=3960 $Y=-6860
X22 6 M2_M1_CDNS_765070438335 $T=4210 -5370 0 0 $X=3960 $Y=-5500
X23 2 M2_M1_CDNS_765070438335 $T=4540 -5740 0 0 $X=4290 $Y=-5870
X24 7 M2_M1_CDNS_765070438335 $T=4960 -4960 0 0 $X=4710 $Y=-5090
X25 7 M2_M1_CDNS_765070438335 $T=4960 -2500 0 0 $X=4710 $Y=-2630
X26 3 M1_PO_CDNS_765070438336 $T=3500 -4810 0 0 $X=3260 $Y=-4910
X27 6 M1_PO_CDNS_765070438336 $T=4210 -6730 0 0 $X=3970 $Y=-6830
X28 6 M1_PO_CDNS_765070438336 $T=4210 -5370 0 0 $X=3970 $Y=-5470
X29 2 M1_PO_CDNS_765070438336 $T=4540 -5740 0 0 $X=4300 $Y=-5840
X30 7 M1_PO_CDNS_765070438336 $T=4960 -4960 0 0 $X=4720 $Y=-5060
X31 7 M1_PO_CDNS_765070438336 $T=4960 -2500 0 0 $X=4720 $Y=-2600
X32 8 2 3 9 pmos1v_CDNS_765070438330 $T=5520 -3500 0 270 $X=5320 $Y=-4010
X33 8 6 7 9 pmos1v_CDNS_765070438330 $T=5520 -2570 0 270 $X=5320 $Y=-3080
X34 5 7 4 9 8 pmos1v_CDNS_765070438331 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X35 9 6 10 nmos1v_CDNS_765070438332 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X36 4 8 6 9 pmos1v_CDNS_765070438333 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X37 8 2 11 9 pmos1v_CDNS_765070438334 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X38 10 6 11 9 8 pmos1v_CDNS_765070438335 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X39 9 10 2 9 nmos1v_CDNS_765070438336 $T=1570 -6390 0 270 $X=1370 $Y=-6840
X40 1 5 2 9 nmos1v_CDNS_765070438336 $T=1570 -4430 0 270 $X=1370 $Y=-4880
X41 1 6 9 nmos1v_CDNS_765070438337 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X42 3 5 12 9 nmos1v_CDNS_765070438338 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X43 9 7 12 nmos1v_CDNS_765070438339 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X44 4 2 8 9 pmos1v_CDNS_7650704383310 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X45 4 3 5 9 8 pmos1v_CDNS_7650704383311 $T=5520 -4430 0 270 $X=5320 $Y=-4760
X46 9 2 3 nmos1v_CDNS_7650704383312 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X47 9 6 7 nmos1v_CDNS_7650704383312 $T=1580 -2570 0 270 $X=1020 $Y=-3080
M0 9 2 10 9 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 1 2 5 9 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M2 8 3 2 8 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.455 scb=0.0418535 scc=0.0112996 $X=5520 $Y=-3590 $dt=1
M3 8 7 6 8 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=5520 $Y=-2660 $dt=1
.ends HAdder
