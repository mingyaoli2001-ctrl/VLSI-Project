* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : MAC                                          *
* Netlisted  : Sat Dec 13 12:39:58 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593021                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593021 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593021

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR a vdd gnd f b 6 7
*.DEVICECLIMB
** N=7 EP=7 FDC=4
X20 gnd gnd a 6 nmos1v_CDNS_765647593021 $T=420 800 0 0 $X=0 $Y=240
X21 f gnd b 6 nmos1v_CDNS_765647593021 $T=1440 800 1 180 $X=930 $Y=240
X22 f gnd 7 a nmos1v_CDNS_765647593021 $T=2280 800 0 0 $X=1860 $Y=240
X23 gnd gnd b 7 nmos1v_CDNS_765647593021 $T=3300 800 1 180 $X=2790 $Y=240
.ends XOR

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593022                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593022 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=6.70537 scb=0.00332581 scc=2.28218e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593022

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593024                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593024 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593024

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593027                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593027 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.78406 scb=0.00345708 scc=2.49632e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593027

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND b a Vdd gnd Vout 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X7 gnd Vout 6 nmos1v_CDNS_765647593022 $T=4560 -2770 0 0 $X=3980 $Y=-2970
X9 gnd b 7 nmos1v_CDNS_765647593024 $T=2230 -2760 1 180 $X=1940 $Y=-2960
X12 6 a 7 gnd nmos1v_CDNS_765647593027 $T=2020 -2760 1 180 $X=1510 $Y=-2960
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_765647593028                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_765647593028 1 2 3 4
** N=5 EP=4 FDC=1
M0 4 3 1 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_765647593028

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_765647593029                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_765647593029 1 2 3 4
** N=4 EP=4 FDC=1
M0 4 3 1 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_765647593029

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CLA_logic                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CLA_logic p1 g1 c0 vdd gnd p2 g2 cout1 p3 g3
+ cout2 p4 cout3 g4 cout4 19 29
*.DEVICECLIMB
** N=39 EP=17 FDC=54
X109 gnd gnd p1 30 nmos1v_CDNS_765647593021 $T=1030 800 0 0 $X=610 $Y=240
X110 30 gnd c0 16 nmos1v_CDNS_765647593021 $T=1960 800 0 0 $X=1540 $Y=240
X111 gnd gnd p2 31 nmos1v_CDNS_765647593021 $T=4750 800 0 0 $X=4330 $Y=240
X112 31 gnd g1 17 nmos1v_CDNS_765647593021 $T=7540 800 0 0 $X=7120 $Y=240
X113 gnd gnd g2 17 nmos1v_CDNS_765647593021 $T=8560 800 1 180 $X=8050 $Y=240
X114 gnd gnd 17 cout2 nmos1v_CDNS_765647593021 $T=9400 800 0 0 $X=8980 $Y=240
X115 32 gnd p1 33 nmos1v_CDNS_765647593021 $T=12190 800 0 0 $X=11770 $Y=240
X116 33 gnd c0 18 nmos1v_CDNS_765647593021 $T=13120 800 0 0 $X=12700 $Y=240
X117 34 gnd g2 18 nmos1v_CDNS_765647593021 $T=14980 800 0 0 $X=14560 $Y=240
X118 gnd gnd g3 18 nmos1v_CDNS_765647593021 $T=16000 800 1 180 $X=15490 $Y=240
X119 gnd gnd 18 cout3 nmos1v_CDNS_765647593021 $T=16840 800 0 0 $X=16420 $Y=240
X120 35 gnd p3 36 nmos1v_CDNS_765647593021 $T=18700 800 0 0 $X=18280 $Y=240
X121 36 gnd g2 19 nmos1v_CDNS_765647593021 $T=23350 800 0 0 $X=22930 $Y=240
X122 gnd gnd 19 cout4 nmos1v_CDNS_765647593021 $T=26140 800 0 0 $X=25720 $Y=240
X326 vdd vdd p1 16 pmos1v_CDNS_765647593028 $T=1030 8610 1 0 $X=610 $Y=8170
X327 20 vdd c0 16 pmos1v_CDNS_765647593028 $T=2050 8610 0 180 $X=1540 $Y=8170
X328 22 vdd p1 17 pmos1v_CDNS_765647593028 $T=5770 8610 0 180 $X=5260 $Y=8170
X329 vdd vdd 18 cout3 pmos1v_CDNS_765647593028 $T=16840 8610 1 0 $X=16420 $Y=8170
X330 29 vdd p3 19 pmos1v_CDNS_765647593028 $T=18790 8610 0 180 $X=18280 $Y=8170
X331 28 vdd c0 19 pmos1v_CDNS_765647593028 $T=21580 8610 0 180 $X=21070 $Y=8170
X332 29 vdd g3 26 pmos1v_CDNS_765647593028 $T=24370 8610 0 180 $X=23860 $Y=8170
X333 gnd gnd g1 16 nmos1v_CDNS_765647593029 $T=2980 1040 0 180 $X=2470 $Y=240
X334 gnd gnd 16 cout1 nmos1v_CDNS_765647593029 $T=3820 1040 1 0 $X=3400 $Y=240
X335 31 gnd p1 37 nmos1v_CDNS_765647593029 $T=5680 1040 1 0 $X=5260 $Y=240
X336 37 gnd c0 17 nmos1v_CDNS_765647593029 $T=6610 1040 1 0 $X=6190 $Y=240
X337 gnd gnd p3 34 nmos1v_CDNS_765647593029 $T=10330 1040 1 0 $X=9910 $Y=240
X338 34 gnd p2 32 nmos1v_CDNS_765647593029 $T=11260 1040 1 0 $X=10840 $Y=240
X339 32 gnd g1 18 nmos1v_CDNS_765647593029 $T=14050 1040 1 0 $X=13630 $Y=240
X340 gnd gnd p4 35 nmos1v_CDNS_765647593029 $T=17770 1040 1 0 $X=17350 $Y=240
X341 36 gnd p2 38 nmos1v_CDNS_765647593029 $T=19630 1040 1 0 $X=19210 $Y=240
X342 38 gnd p1 39 nmos1v_CDNS_765647593029 $T=20560 1040 1 0 $X=20140 $Y=240
X343 39 gnd c0 19 nmos1v_CDNS_765647593029 $T=21490 1040 1 0 $X=21070 $Y=240
X344 38 gnd g1 19 nmos1v_CDNS_765647593029 $T=22420 1040 1 0 $X=22000 $Y=240
X345 35 gnd g3 19 nmos1v_CDNS_765647593029 $T=24280 1040 1 0 $X=23860 $Y=240
X346 gnd gnd g4 19 nmos1v_CDNS_765647593029 $T=25300 1040 0 180 $X=24790 $Y=240
M0 vdd g1 20 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=2890 $Y=8370 $dt=1
M1 cout1 16 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=3820 $Y=8370 $dt=1
M2 17 p2 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=4750 $Y=8370 $dt=1
M3 21 c0 17 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=6610 $Y=8370 $dt=1
M4 22 g1 21 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=7540 $Y=8370 $dt=1
M5 vdd g2 22 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=8470 $Y=8370 $dt=1
M6 cout2 17 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=9400 $Y=8370 $dt=1
M7 18 p3 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=10330 $Y=8370 $dt=1
M8 23 p2 18 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=11260 $Y=8370 $dt=1
M9 24 p1 18 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=12190 $Y=8370 $dt=1
M10 25 c0 18 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=13120 $Y=8370 $dt=1
M11 24 g1 25 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14050 $Y=8370 $dt=1
M12 23 g2 24 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=14980 $Y=8370 $dt=1
M13 vdd g3 23 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=15910 $Y=8370 $dt=1
M14 19 p4 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=17770 $Y=8370 $dt=1
M15 26 p2 19 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=19630 $Y=8370 $dt=1
M16 27 p1 19 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=20560 $Y=8370 $dt=1
M17 27 g1 28 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=22420 $Y=8370 $dt=1
M18 26 g2 27 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=23350 $Y=8370 $dt=1
.ends 4bit_CLA_logic

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930210                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930210 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930210

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930211                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930211 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930211

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930212                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930212 1 2 3
** N=4 EP=3 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930212

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930213                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930213 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930213

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930214                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930214 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930214

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930216                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930216 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930216

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930217                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930217 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930217

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7656475930218                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7656475930218 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7656475930218

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930219                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930219 1 2 3
** N=4 EP=3 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=6.86517 scb=0.00359333 scc=2.73027e-05 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930219

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7656475930220                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7656475930220 1 2 3 5
** N=5 EP=4 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=78.5337 scb=0.0310796 scc=0.00873963 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7656475930220

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder sum gnd carry a b vdd
** N=12 EP=6 FDC=16
X19 gnd gnd a 8 nmos1v_CDNS_765647593021 $T=1570 -3500 0 270 $X=1010 $Y=-4010
X20 gnd gnd b 7 nmos1v_CDNS_765647593021 $T=1580 -2570 0 270 $X=1020 $Y=-3080
X36 sum b 9 vdd pmos1v_CDNS_7656475930210 $T=5520 -4930 1 90 $X=5320 $Y=-5170
X37 gnd 7 carry nmos1v_CDNS_7656475930211 $T=1570 -6890 1 90 $X=1370 $Y=-7310
X38 9 vdd 7 pmos1v_CDNS_7656475930212 $T=5520 -5340 1 90 $X=5320 $Y=-5700
X39 vdd 8 11 pmos1v_CDNS_7656475930213 $T=5520 -6590 0 270 $X=5320 $Y=-6880
X40 carry 7 11 vdd pmos1v_CDNS_7656475930214 $T=5520 -6800 0 270 $X=5320 $Y=-7310
X43 10 7 gnd nmos1v_CDNS_7656475930216 $T=1570 -5460 0 270 $X=1370 $Y=-5970
X44 a sum 12 gnd nmos1v_CDNS_7656475930217 $T=1570 -4930 1 90 $X=1370 $Y=-5130
X45 gnd b 12 nmos1v_CDNS_7656475930218 $T=1570 -5140 1 90 $X=1370 $Y=-5500
X46 9 8 vdd pmos1v_CDNS_7656475930219 $T=5520 -5660 0 270 $X=5320 $Y=-6170
X47 9 a sum vdd pmos1v_CDNS_7656475930220 $T=5520 -4430 0 270 $X=5320 $Y=-4760
M0 gnd 8 carry gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6480 $dt=0
M1 10 8 sum gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4520 $dt=0
M2 vdd a 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=100.171 scb=0.0396101 scc=0.0112296 $X=5520 $Y=-3590 $dt=1
M3 vdd b 7 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=118.462 scb=0.0629606 scc=0.0138757 $X=5520 $Y=-2660 $dt=1
.ends HAdder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MAC                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MAC c<0> c<10> c<11> c<12> c<13> c<14> c<15> c<1> c<2> c<3>
+ c<4> c<5> c<6> c<7> c<8> c<9> gnd mac<0> mac<10> mac<11>
+ mac<12> mac<13> mac<14> mac<15> mac<16> mac<1> mac<2> mac<3> mac<4> mac<5>
+ mac<6> mac<7> mac<8> mac<9> s<0> s<10> s<11> s<12> s<13> s<14>
+ s<15> s<1> s<2> s<3> s<4> s<5> s<6> s<7> s<8> s<9>
+ vdd
** N=291 EP=51 FDC=570
X181 17 vdd gnd mac<9> 1 163 100 XOR $T=640 25900 1 0 $X=640 $Y=21200
X182 s<8> vdd gnd 2 c<8> 164 101 XOR $T=4740 40010 1 0 $X=4740 $Y=35310
X183 18 vdd gnd mac<8> 2 165 102 XOR $T=9740 25900 0 180 $X=6020 $Y=21200
X184 19 vdd gnd mac<15> 4 166 103 XOR $T=17180 4700 0 180 $X=13460 $Y=0
X185 20 vdd gnd mac<7> 5 167 104 XOR $T=17180 25900 0 180 $X=13460 $Y=21200
X186 s<15> vdd gnd 4 c<15> 168 105 XOR $T=13530 18810 1 0 $X=13530 $Y=14110
X187 s<7> vdd gnd 5 c<7> 169 106 XOR $T=13530 40010 1 0 $X=13530 $Y=35310
X188 21 vdd gnd mac<14> 6 170 107 XOR $T=22760 4700 0 180 $X=19040 $Y=0
X189 22 vdd gnd mac<6> 7 171 108 XOR $T=22760 25900 0 180 $X=19040 $Y=21200
X190 s<14> vdd gnd 6 c<14> 172 109 XOR $T=19120 18810 1 0 $X=19120 $Y=14110
X191 s<6> vdd gnd 7 c<6> 173 110 XOR $T=19120 40010 1 0 $X=19120 $Y=35310
X192 23 vdd gnd mac<13> 8 174 111 XOR $T=26810 4700 0 180 $X=23090 $Y=0
X193 24 vdd gnd mac<5> 9 175 112 XOR $T=26810 25900 0 180 $X=23090 $Y=21200
X194 s<13> vdd gnd 8 c<13> 176 113 XOR $T=31140 18810 0 180 $X=27420 $Y=14110
X195 s<5> vdd gnd 9 c<5> 177 114 XOR $T=31140 40010 0 180 $X=27420 $Y=35310
X196 s<12> vdd gnd 10 c<12> 178 115 XOR $T=31430 18810 1 0 $X=31430 $Y=14110
X197 s<4> vdd gnd 11 c<4> 179 116 XOR $T=31430 40010 1 0 $X=31430 $Y=35310
X198 25 vdd gnd mac<12> 10 180 117 XOR $T=36470 4700 0 180 $X=32750 $Y=0
X199 26 vdd gnd mac<4> 11 181 118 XOR $T=36470 25900 0 180 $X=32750 $Y=21200
X200 27 vdd gnd mac<11> 12 182 119 XOR $T=43890 4700 0 180 $X=40170 $Y=0
X201 28 vdd gnd mac<3> 13 183 120 XOR $T=43890 25900 0 180 $X=40170 $Y=21200
X202 s<11> vdd gnd 12 c<11> 184 121 XOR $T=40220 18810 1 0 $X=40220 $Y=14110
X203 s<3> vdd gnd 13 c<3> 185 122 XOR $T=40220 40010 1 0 $X=40220 $Y=35310
X204 29 vdd gnd mac<10> 14 186 123 XOR $T=49450 4700 0 180 $X=45730 $Y=0
X205 30 vdd gnd mac<2> 15 187 124 XOR $T=49450 25900 0 180 $X=45730 $Y=21200
X206 s<10> vdd gnd 14 c<10> 188 125 XOR $T=45810 18810 1 0 $X=45810 $Y=14110
X207 s<2> vdd gnd 15 c<2> 189 126 XOR $T=45810 40010 1 0 $X=45810 $Y=35310
X208 90 vdd gnd mac<1> 16 190 127 XOR $T=49650 25900 1 0 $X=49650 $Y=21200
X209 s<9> vdd gnd 1 c<9> 191 128 XOR $T=57790 18810 0 180 $X=54070 $Y=14110
X210 s<1> vdd gnd 16 c<1> 192 129 XOR $T=57790 40010 0 180 $X=54070 $Y=35310
X211 c<8> s<8> vdd gnd 31 130 AND $T=3670 43110 0 0 $X=4740 $Y=40010
X212 c<15> s<15> vdd gnd 32 131 AND $T=12460 21910 0 0 $X=13530 $Y=18810
X213 c<7> s<7> vdd gnd 33 132 AND $T=12460 43110 0 0 $X=13530 $Y=40010
X214 c<14> s<14> vdd gnd 34 133 AND $T=18050 21910 0 0 $X=19120 $Y=18810
X215 c<6> s<6> vdd gnd 35 134 AND $T=18050 43110 0 0 $X=19120 $Y=40010
X216 c<13> s<13> vdd gnd 36 135 AND $T=32170 21910 1 180 $X=26920 $Y=18810
X217 c<5> s<5> vdd gnd 37 136 AND $T=32170 43110 1 180 $X=26920 $Y=40010
X218 c<12> s<12> vdd gnd 38 137 AND $T=30360 21910 0 0 $X=31430 $Y=18810
X219 c<4> s<4> vdd gnd 39 138 AND $T=30360 43110 0 0 $X=31430 $Y=40010
X220 c<11> s<11> vdd gnd 40 139 AND $T=39150 21910 0 0 $X=40220 $Y=18810
X221 c<3> s<3> vdd gnd 41 140 AND $T=39150 43110 0 0 $X=40220 $Y=40010
X222 c<10> s<10> vdd gnd 42 141 AND $T=44740 21910 0 0 $X=45810 $Y=18810
X223 c<2> s<2> vdd gnd 43 142 AND $T=44740 43110 0 0 $X=45810 $Y=40010
X224 c<9> s<9> vdd gnd 44 143 AND $T=58860 21910 1 180 $X=53610 $Y=18810
X225 c<1> s<1> vdd gnd 45 144 AND $T=58860 43110 1 180 $X=53610 $Y=40010
X226 8 36 23 vdd gnd 6 34 21 4 32
+ 19 94 mac<16> 95 96 148 256 4bit_CLA_logic $T=26970 4700 1 180 $X=320 $Y=4700
X227 9 37 24 vdd gnd 7 35 22 5 33
+ 20 2 18 31 17 152 266 4bit_CLA_logic $T=26970 25900 1 180 $X=320 $Y=25900
X228 1 44 17 vdd gnd 14 42 29 12 40
+ 27 10 25 38 23 156 276 4bit_CLA_logic $T=53660 4700 1 180 $X=27010 $Y=4700
X229 16 45 90 vdd gnd 15 43 30 13 41
+ 28 11 26 39 24 160 286 4bit_CLA_logic $T=53660 25900 1 180 $X=27010 $Y=25900
X230 mac<0> gnd 90 s<0> c<0> vdd HAdder $T=62720 27380 1 90 $X=53760 $Y=28180
M0 vdd 148 96 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=13070 $dt=1
M1 vdd 152 17 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=23.1856 scb=0.0241633 scc=0.00264686 $X=740 $Y=34270 $dt=1
M2 163 17 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=1060 $Y=22000 $dt=1
M3 256 95 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=13070 $dt=1
M4 266 31 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=4.89541 scb=0.000812888 scc=7.58777e-07 $X=1670 $Y=34270 $dt=1
M5 mac<9> 1 17 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=1990 $Y=22000 $dt=1
M6 163 100 mac<9> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=2920 $Y=22000 $dt=1
M7 vdd 1 100 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=3850 $Y=22000 $dt=1
M8 164 s<8> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=5160 $Y=36110 $dt=1
M9 130 s<8> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=5600 $Y=41790 $dt=1
M10 vdd c<8> 130 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=6010 $Y=41790 $dt=1
M11 2 c<8> s<8> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=6090 $Y=36110 $dt=1
M12 102 2 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=6440 $Y=22000 $dt=1
M13 164 101 2 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7020 $Y=36110 $dt=1
M14 mac<8> 102 165 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=7370 $Y=22000 $dt=1
M15 vdd c<8> 101 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=7950 $Y=36110 $dt=1
M16 31 130 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=8230 $Y=41600 $dt=1
M17 18 2 mac<8> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=8300 $Y=22000 $dt=1
M18 vdd 18 165 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=9230 $Y=22000 $dt=1
M19 103 4 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=13880 $Y=800 $dt=1
M20 104 5 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=115.144 scb=0.0588049 scc=0.0138331 $X=13880 $Y=22000 $dt=1
M21 168 s<15> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=14910 $dt=1
M22 169 s<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=13950 $Y=36110 $dt=1
M23 131 s<15> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=30.29 scb=0.029437 scc=0.00332952 $X=14390 $Y=20590 $dt=1
M24 132 s<7> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=14390 $Y=41790 $dt=1
M25 vdd c<15> 131 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=28.0435 scb=0.0261338 scc=0.00329543 $X=14800 $Y=20590 $dt=1
M26 vdd c<7> 132 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=14800 $Y=41790 $dt=1
M27 mac<15> 103 166 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=14810 $Y=800 $dt=1
M28 mac<7> 104 167 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=96.854 scb=0.0354545 scc=0.011187 $X=14810 $Y=22000 $dt=1
M29 4 c<15> s<15> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=14910 $dt=1
M30 5 c<7> s<7> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=14880 $Y=36110 $dt=1
M31 19 4 mac<15> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=15740 $Y=800 $dt=1
M32 20 5 mac<7> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=15740 $Y=22000 $dt=1
M33 168 105 4 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=14910 $dt=1
M34 169 106 5 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=15810 $Y=36110 $dt=1
M35 vdd 19 166 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=16670 $Y=800 $dt=1
M36 vdd 20 167 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=16670 $Y=22000 $dt=1
M37 vdd c<15> 105 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=14910 $dt=1
M38 vdd c<7> 106 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=16740 $Y=36110 $dt=1
M39 32 131 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=17020 $Y=20400 $dt=1
M40 33 132 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=17020 $Y=41600 $dt=1
M41 107 6 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=19460 $Y=800 $dt=1
M42 108 7 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=19460 $Y=22000 $dt=1
M43 172 s<14> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=14910 $dt=1
M44 173 s<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=19540 $Y=36110 $dt=1
M45 133 s<14> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=19980 $Y=20590 $dt=1
M46 134 s<6> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=19980 $Y=41790 $dt=1
M47 mac<14> 107 170 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=20390 $Y=800 $dt=1
M48 vdd c<14> 133 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=20390 $Y=20590 $dt=1
M49 mac<6> 108 171 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=20390 $Y=22000 $dt=1
M50 vdd c<6> 134 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=20390 $Y=41790 $dt=1
M51 6 c<14> s<14> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=14910 $dt=1
M52 7 c<6> s<6> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=20470 $Y=36110 $dt=1
M53 21 6 mac<14> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=21320 $Y=800 $dt=1
M54 22 7 mac<6> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=21320 $Y=22000 $dt=1
M55 172 109 6 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=14910 $dt=1
M56 173 110 7 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=21400 $Y=36110 $dt=1
M57 vdd 21 170 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=22250 $Y=800 $dt=1
M58 vdd 22 171 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=22250 $Y=22000 $dt=1
M59 vdd c<14> 109 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=14910 $dt=1
M60 vdd c<6> 110 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=22330 $Y=36110 $dt=1
M61 34 133 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=22610 $Y=20400 $dt=1
M62 35 134 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=22610 $Y=41600 $dt=1
M63 111 8 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=23510 $Y=800 $dt=1
M64 112 9 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=23510 $Y=22000 $dt=1
M65 mac<13> 111 174 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=101.24 scb=0.0428046 scc=0.0113759 $X=24440 $Y=800 $dt=1
M66 mac<5> 112 175 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=24440 $Y=22000 $dt=1
M67 23 8 mac<13> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=25370 $Y=800 $dt=1
M68 24 9 mac<5> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=25370 $Y=22000 $dt=1
M69 vdd 23 174 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=26300 $Y=800 $dt=1
M70 vdd 24 175 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=26300 $Y=22000 $dt=1
M71 vdd 156 23 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=13070 $dt=1
M72 vdd 160 24 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=27430 $Y=34270 $dt=1
M73 vdd 135 36 vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=27520 $Y=20400 $dt=1
M74 vdd 136 37 vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=27520 $Y=41600 $dt=1
M75 113 c<13> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=14910 $dt=1
M76 114 c<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=27840 $Y=36110 $dt=1
M77 276 38 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=13070 $dt=1
M78 286 39 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.73438 scb=0.00013556 scc=4.76679e-09 $X=28360 $Y=34270 $dt=1
M79 8 113 176 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=14910 $dt=1
M80 9 114 177 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=28770 $Y=36110 $dt=1
M81 s<13> c<13> 8 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=14910 $dt=1
M82 s<5> c<5> 9 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=29700 $Y=36110 $dt=1
M83 135 c<13> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=29740 $Y=20590 $dt=1
M84 136 c<5> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=29740 $Y=41790 $dt=1
M85 vdd s<13> 135 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=30150 $Y=20590 $dt=1
M86 vdd s<5> 136 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=30150 $Y=41790 $dt=1
M87 vdd s<13> 176 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=14910 $dt=1
M88 vdd s<5> 177 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=30630 $Y=36110 $dt=1
M89 178 s<12> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=14910 $dt=1
M90 179 s<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=31850 $Y=36110 $dt=1
M91 137 s<12> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32290 $Y=20590 $dt=1
M92 138 s<4> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32290 $Y=41790 $dt=1
M93 vdd c<12> 137 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=32700 $Y=20590 $dt=1
M94 vdd c<4> 138 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=43.0969 scb=0.0465601 scc=0.00538363 $X=32700 $Y=41790 $dt=1
M95 10 c<12> s<12> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=14910 $dt=1
M96 11 c<4> s<4> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=32780 $Y=36110 $dt=1
M97 117 10 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=33170 $Y=800 $dt=1
M98 118 11 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=33170 $Y=22000 $dt=1
M99 178 115 10 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=14910 $dt=1
M100 179 116 11 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=33710 $Y=36110 $dt=1
M101 mac<12> 117 180 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=34100 $Y=800 $dt=1
M102 mac<4> 118 181 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=34100 $Y=22000 $dt=1
M103 vdd c<12> 115 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=14910 $dt=1
M104 vdd c<4> 116 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=34640 $Y=36110 $dt=1
M105 38 137 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=34920 $Y=20400 $dt=1
M106 39 138 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=34920 $Y=41600 $dt=1
M107 25 10 mac<12> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=35030 $Y=800 $dt=1
M108 26 11 mac<4> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35030 $Y=22000 $dt=1
M109 vdd 25 180 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=35960 $Y=800 $dt=1
M110 vdd 26 181 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=35960 $Y=22000 $dt=1
M111 119 12 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=40590 $Y=800 $dt=1
M112 120 13 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=40590 $Y=22000 $dt=1
M113 184 s<11> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=14910 $dt=1
M114 185 s<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=40640 $Y=36110 $dt=1
M115 139 s<11> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41080 $Y=20590 $dt=1
M116 140 s<3> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=41080 $Y=41790 $dt=1
M117 vdd c<11> 139 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=41490 $Y=20590 $dt=1
M118 vdd c<3> 140 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=41490 $Y=41790 $dt=1
M119 mac<11> 119 182 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=41520 $Y=800 $dt=1
M120 mac<3> 120 183 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=41520 $Y=22000 $dt=1
M121 12 c<11> s<11> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=14910 $dt=1
M122 13 c<3> s<3> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=41570 $Y=36110 $dt=1
M123 27 12 mac<11> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=42450 $Y=800 $dt=1
M124 28 13 mac<3> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=42450 $Y=22000 $dt=1
M125 184 121 12 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=14910 $dt=1
M126 185 122 13 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=42500 $Y=36110 $dt=1
M127 vdd 27 182 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=43380 $Y=800 $dt=1
M128 vdd 28 183 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=43380 $Y=22000 $dt=1
M129 vdd c<11> 121 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=14910 $dt=1
M130 vdd c<3> 122 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=43430 $Y=36110 $dt=1
M131 40 139 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=43710 $Y=20400 $dt=1
M132 41 140 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=43710 $Y=41600 $dt=1
M133 123 14 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=46150 $Y=800 $dt=1
M134 124 15 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=46150 $Y=22000 $dt=1
M135 188 s<10> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=14910 $dt=1
M136 189 s<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=46230 $Y=36110 $dt=1
M137 141 s<10> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=46670 $Y=20590 $dt=1
M138 142 s<2> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=46670 $Y=41790 $dt=1
M139 mac<10> 123 186 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=47080 $Y=800 $dt=1
M140 vdd c<10> 141 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=26.8513 scb=0.0254253 scc=0.00329461 $X=47080 $Y=20590 $dt=1
M141 mac<2> 124 187 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=47080 $Y=22000 $dt=1
M142 vdd c<2> 142 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=47080 $Y=41790 $dt=1
M143 14 c<10> s<10> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=14910 $dt=1
M144 15 c<2> s<2> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=47160 $Y=36110 $dt=1
M145 29 14 mac<10> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=102.402 scb=0.043482 scc=0.0113766 $X=48010 $Y=800 $dt=1
M146 30 15 mac<2> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48010 $Y=22000 $dt=1
M147 188 125 14 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=14910 $dt=1
M148 189 126 15 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=48090 $Y=36110 $dt=1
M149 vdd 29 186 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=48940 $Y=800 $dt=1
M150 vdd 30 187 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=48940 $Y=22000 $dt=1
M151 vdd c<10> 125 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=14910 $dt=1
M152 vdd c<2> 126 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=49020 $Y=36110 $dt=1
M153 42 141 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=49300 $Y=20400 $dt=1
M154 43 142 vdd vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=49300 $Y=41600 $dt=1
M155 190 90 vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=50070 $Y=22000 $dt=1
M156 mac<1> 16 90 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51000 $Y=22000 $dt=1
M157 190 127 mac<1> vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=51930 $Y=22000 $dt=1
M158 vdd 16 127 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.693 scb=0.0347772 scc=0.0111862 $X=52860 $Y=22000 $dt=1
M159 vdd 143 44 vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=58.8484 scb=0.0285532 scc=0.00672169 $X=54210 $Y=20400 $dt=1
M160 vdd 144 45 vdd g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=93.2539 scb=0.0709721 scc=0.0112581 $X=54210 $Y=41600 $dt=1
M161 128 c<9> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=14910 $dt=1
M162 129 c<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=54490 $Y=36110 $dt=1
M163 1 128 191 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=14910 $dt=1
M164 16 129 192 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.3993 scb=0.0347075 scc=0.0111862 $X=55420 $Y=36110 $dt=1
M165 s<9> c<9> 1 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=14910 $dt=1
M166 s<1> c<1> 16 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=95.6441 scb=0.0347702 scc=0.0111862 $X=56350 $Y=36110 $dt=1
M167 143 c<9> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=29.0043 scb=0.0273456 scc=0.00330147 $X=56430 $Y=20590 $dt=1
M168 144 c<1> vdd vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=45.2499 scb=0.0484803 scc=0.00539049 $X=56430 $Y=41790 $dt=1
M169 vdd s<9> 143 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=33.5338 scb=0.0350848 scc=0.00355838 $X=56840 $Y=20590 $dt=1
M170 vdd s<1> 144 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=49.7794 scb=0.0562196 scc=0.00564739 $X=56840 $Y=41790 $dt=1
M171 vdd s<9> 191 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=14910 $dt=1
M172 vdd s<1> 192 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=99.4486 scb=0.0397911 scc=0.0112458 $X=57280 $Y=36110 $dt=1
.ends MAC
