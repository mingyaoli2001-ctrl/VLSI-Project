* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : HAdder                                       *
* Netlisted  : Fri Dec  5 01:26:36 2025                     *
* PVS Version: 23.11-s036 Wed Jan 17 18:11:41 PST 2024      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764915992331                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764915992331 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764915992331

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764915992332                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764915992332 1 2 3
** N=4 EP=3 FDC=1
M0 1 3 2 2 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=5.5e-07 sca=96.8699 scb=0.035625 scc=0.0111877 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764915992332

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764915992333                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764915992333 1 2 3 5
** N=5 EP=4 FDC=1
M0 3 2 1 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=7.55e-07 sca=96.8213 scb=0.0356156 scc=0.0111877 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764915992333

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764915992334                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764915992334 1 2 3
** N=4 EP=3 FDC=1
M0 3 2 1 1 g45p1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=105.232 scb=0.0480039 scc=0.0116671 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764915992334

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_764915992335                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_764915992335 1 2 3 5
** N=5 EP=4 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=116.273 scb=0.0596433 scc=0.0138346 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_764915992335

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764915992337                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764915992337 1 2 3
** N=3 EP=3 FDC=1
M0 1 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764915992337

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764915992338                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764915992338 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 1 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=7.2e-15 PD=5.6e-07 PS=3.6e-07 fw=1.2e-07 sa=4.5e-07 sb=3.45e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764915992338

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_764915992339                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_764915992339 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.92e-14 PD=3.6e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=4.5e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_764915992339

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7649159923310                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7649159923310 1 2 3
** N=4 EP=3 FDC=1
M0 1 2 3 3 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=7.55e-07 sb=1.4e-07 sca=97.4578 scb=0.0358666 scc=0.0111878 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7649159923310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_7649159923311                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_7649159923311 1 2 3 5
** N=5 EP=4 FDC=1
M0 2 1 3 5 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.92e-14 PD=5.6e-07 PS=5.6e-07 fw=1.2e-07 sa=5.5e-07 sb=3.45e-07 sca=96.8213 scb=0.0356156 scc=0.0111877 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_7649159923311

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7649159923312                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7649159923312 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7649159923312

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAdder                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAdder a b carry gnd sum vdd
** N=12 EP=6 FDC=16
X23 gnd 10 carry nmos1v_CDNS_764915992331 $T=1570 -6910 1 90 $X=1370 $Y=-7330
X24 7 vdd 10 pmos1v_CDNS_764915992332 $T=5040 -5340 1 90 $X=4840 $Y=-5700
X25 7 a sum vdd pmos1v_CDNS_764915992333 $T=5040 -4430 0 270 $X=4840 $Y=-4880
X26 vdd 1 11 pmos1v_CDNS_764915992334 $T=5040 -6590 0 270 $X=4840 $Y=-6880
X27 carry 10 11 vdd pmos1v_CDNS_764915992335 $T=5040 -6800 0 270 $X=4840 $Y=-7310
X30 5 10 gnd nmos1v_CDNS_764915992337 $T=1570 -5480 0 270 $X=1370 $Y=-5990
X31 a sum 12 gnd nmos1v_CDNS_764915992338 $T=1570 -4950 1 90 $X=1370 $Y=-5150
X32 gnd b 12 nmos1v_CDNS_764915992339 $T=1570 -5160 1 90 $X=1370 $Y=-5520
X33 7 1 vdd pmos1v_CDNS_7649159923310 $T=5040 -5660 0 270 $X=4840 $Y=-6170
X34 b sum 7 vdd pmos1v_CDNS_7649159923311 $T=5040 -4930 1 90 $X=4840 $Y=-5170
X35 gnd 1 a nmos1v_CDNS_7649159923312 $T=1570 -3520 0 270 $X=1010 $Y=-4030
X36 gnd 10 b nmos1v_CDNS_7649159923312 $T=1580 -2590 0 270 $X=1020 $Y=-3100
M0 gnd 1 carry gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-6500 $dt=0
M1 5 1 sum gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=6.55e-07 sb=1.4e-07 sca=3.69959 scb=0.00013007 scc=4.39142e-09 $X=1570 $Y=-4540 $dt=0
M2 vdd a 1 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=97.9823 scb=0.0362929 scc=0.0111885 $X=5040 $Y=-3590 $dt=1
M3 vdd b 10 vdd g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=120.692 scb=0.0668324 scc=0.0140227 $X=5040 $Y=-2660 $dt=1
.ends HAdder
